library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity internalram is
  port (
    CLK:              in std_logic;
    EN:               in std_logic;
    ADDR:             in std_logic_vector(12 downto 2);
    DO:               out std_logic_vector(31 downto 0)
  );
end entity internalram;

architecture behave of internalram is

begin

process(CLK)
variable iaddr: natural;
begin
  if rising_edge(CLK) then
   if EN='1' then
   iaddr := to_integer(unsigned(ADDR));
     case iaddr is 
      when 0 => DO <= x"ffff6000"; 
      when 1 => DO <= x"7fcf8000"; 
      when 2 => DO <= x"70207042"; 
      when 3 => DO <= x"72a11012"; 
      when 4 => DO <= x"74219012"; 
      when 5 => DO <= x"40fc800e"; 
      when 6 => DO <= x"70007001"; 
      when 7 => DO <= x"3e313800"; 
      when 8 => DO <= x"3c113800"; 
      when 9 => DO <= x"85114002"; 
      when 10 => DO <= x"3e113800"; 
      when 11 => DO <= x"30003800"; 
      when 12 => DO <= x"800e7000"; 
      when 13 => DO <= x"7631cc0d"; 
      when 14 => DO <= x"40003800"; 
      when 15 => DO <= x"a0006000"; 
      when 16 => DO <= x"70017002"; 
      when 17 => DO <= x"0c130c24"; 
      when 18 => DO <= x"10225ff1"; 
      when 19 => DO <= x"18520725"; 
      when 20 => DO <= x"c50d4100"; 
      when 21 => DO <= x"38006001"; 
      when 22 => DO <= x"5042cea0"; 
      when 23 => DO <= x"41ff3800"; 
      when 24 => DO <= x"18240742"; 
      when 25 => DO <= x"5ff3c12d"; 
      when 26 => DO <= x"41006003"; 
      when 27 => DO <= x"cf0041ff"; 
      when 28 => DO <= x"5044c92d"; 
      when 29 => DO <= x"40053800"; 
      when 30 => DO <= x"4fe03800"; 
      when 31 => DO <= x"0cdc0c1b"; 
      when 32 => DO <= x"800e7000"; 
      when 33 => DO <= x"7481472d"; 
      when 34 => DO <= x"38000c41"; 
      when 35 => DO <= x"442d3800"; 
      when 36 => DO <= x"800e7000"; 
      when 37 => DO <= x"7611462d"; 
      when 38 => DO <= x"38000c41"; 
      when 39 => DO <= x"432d3800"; 
      when 40 => DO <= x"42603800"; 
      when 41 => DO <= x"0c1b0c27"; 
      when 42 => DO <= x"800e7000"; 
      when 43 => DO <= x"748144ad"; 
      when 44 => DO <= x"38000c71"; 
      when 45 => DO <= x"41ad3800"; 
      when 46 => DO <= x"800e7000"; 
      when 47 => DO <= x"761143ad"; 
      when 48 => DO <= x"38000c51"; 
      when 49 => DO <= x"40ad3800"; 
      when 50 => DO <= x"4fe03800"; 
      when 51 => DO <= x"00000000"; 
      when 52 => DO <= x"0cd50c14"; 
      when 53 => DO <= x"70778941"; 
      when 54 => DO <= x"401c8844"; 
      when 55 => DO <= x"40048411"; 
      when 56 => DO <= x"400f5301"; 
      when 57 => DO <= x"6391d081"; 
      when 58 => DO <= x"4700436d"; 
      when 59 => DO <= x"38006007"; 
      when 60 => DO <= x"ce2041ff"; 
      when 61 => DO <= x"5ff73050"; 
      when 62 => DO <= x"38000c18"; 
      when 63 => DO <= x"1a186001"; 
      when 64 => DO <= x"c0e04200"; 
      when 65 => DO <= x"50180cd6"; 
      when 66 => DO <= x"418d3800"; 
      when 67 => DO <= x"0c6d4ec0"; 
      when 68 => DO <= x"380030d0"; 
      when 69 => DO <= x"38000000"; 
      when 70 => DO <= x"00000000"; 
      when 71 => DO <= x"00000000"; 
      when 72 => DO <= x"00008000"; 
      when 73 => DO <= x"70207002"; 
      when 74 => DO <= x"98324004"; 
      when 75 => DO <= x"84334002"; 
      when 76 => DO <= x"6003cf20"; 
      when 77 => DO <= x"41ff3800"; 
      when 78 => DO <= x"101230d0"; 
      when 79 => DO <= x"38007021"; 
      when 80 => DO <= x"24413800"; 
      when 81 => DO <= x"38003800"; 
      when 82 => DO <= x"20413800"; 
      when 83 => DO <= x"84124002"; 
      when 84 => DO <= x"6002cf20"; 
      when 85 => DO <= x"41ff3800"; 
      when 86 => DO <= x"30d03800"; 
      when 87 => DO <= x"70112441"; 
      when 88 => DO <= x"38003800"; 
      when 89 => DO <= x"30d03800"; 
      when 90 => DO <= x"30103800"; 
      when 91 => DO <= x"00000000"; 
      when 92 => DO <= x"00000000"; 
      when 93 => DO <= x"00000000"; 
      when 94 => DO <= x"00008006"; 
      when 95 => DO <= x"7000708d"; 
      when 96 => DO <= x"30d07001"; 
      when 97 => DO <= x"4fe03800"; 
      when 98 => DO <= x"4fe03800"; 
      when 99 => DO <= x"3e5f3800"; 
      when 100 => DO <= x"ffff6000"; 
      when 101 => DO <= x"7fcf180f"; 
      when 102 => DO <= x"101f902f"; 
      when 103 => DO <= x"40fc903f"; 
      when 104 => DO <= x"40f8904f"; 
      when 105 => DO <= x"40f4905f"; 
      when 106 => DO <= x"40f0906f"; 
      when 107 => DO <= x"40ec907f"; 
      when 108 => DO <= x"40e8908f"; 
      when 109 => DO <= x"40e4909f"; 
      when 110 => DO <= x"40e090af"; 
      when 111 => DO <= x"40dc90bf"; 
      when 112 => DO <= x"40d890cf"; 
      when 113 => DO <= x"40d490df"; 
      when 114 => DO <= x"40d090ef"; 
      when 115 => DO <= x"40cc3c51"; 
      when 116 => DO <= x"3800901f"; 
      when 117 => DO <= x"40c83c21"; 
      when 118 => DO <= x"3800901f"; 
      when 119 => DO <= x"40c43c41"; 
      when 120 => DO <= x"3800901f"; 
      when 121 => DO <= x"40c080f1"; 
      when 122 => DO <= x"40c05bcf"; 
      when 123 => DO <= x"c34d4006"; 
      when 124 => DO <= x"3800544f"; 
      when 125 => DO <= x"981f40c0"; 
      when 126 => DO <= x"3e413800"; 
      when 127 => DO <= x"981f40c4"; 
      when 128 => DO <= x"3e213800"; 
      when 129 => DO <= x"981f40c8"; 
      when 130 => DO <= x"3e513800"; 
      when 131 => DO <= x"98ef40cc"; 
      when 132 => DO <= x"98df40d0"; 
      when 133 => DO <= x"98cf40d4"; 
      when 134 => DO <= x"98bf40d8"; 
      when 135 => DO <= x"98af40dc"; 
      when 136 => DO <= x"989f40e0"; 
      when 137 => DO <= x"988f40e4"; 
      when 138 => DO <= x"987f40e8"; 
      when 139 => DO <= x"986f40ec"; 
      when 140 => DO <= x"985f40f0"; 
      when 141 => DO <= x"984f40f4"; 
      when 142 => DO <= x"983f40f8"; 
      when 143 => DO <= x"982f40fc"; 
      when 144 => DO <= x"181f3c5f"; 
      when 145 => DO <= x"38003400"; 
      when 146 => DO <= x"38000c01"; 
      when 147 => DO <= x"0c020c03"; 
      when 148 => DO <= x"0c040c05"; 
      when 149 => DO <= x"0c060c07"; 
      when 150 => DO <= x"0c080c09"; 
      when 151 => DO <= x"0c0a0c0b"; 
      when 152 => DO <= x"30d00c0c"; 
      when 153 => DO <= x"3c113800"; 
      when 154 => DO <= x"30d03800"; 
      when 155 => DO <= x"30d03800"; 
      when 156 => DO <= x"20813800"; 
      when 157 => DO <= x"30d03800"; 
      when 158 => DO <= x"20513800"; 
      when 159 => DO <= x"30d03800"; 
      when 160 => DO <= x"24813800"; 
      when 161 => DO <= x"30d03800"; 
      when 162 => DO <= x"24513800"; 
      when 163 => DO <= x"30d03800"; 
      when 164 => DO <= x"20913800"; 
      when 165 => DO <= x"30d03800"; 
      when 166 => DO <= x"20a13800"; 
      when 167 => DO <= x"30d03800"; 
      when 168 => DO <= x"20b13800"; 
      when 169 => DO <= x"30d03800"; 
      when 170 => DO <= x"20c13800"; 
      when 171 => DO <= x"30d03800"; 
      when 172 => DO <= x"20d13800"; 
      when 173 => DO <= x"30d03800"; 
      when 174 => DO <= x"20e13800"; 
      when 175 => DO <= x"30d03800"; 
      when 176 => DO <= x"24e13800"; 
      when 177 => DO <= x"30d03800"; 
      when 178 => DO <= x"20f13800"; 
      when 179 => DO <= x"30d03800"; 
      when 180 => DO <= x"24613800"; 
      when 181 => DO <= x"30d02071"; 
      when 182 => DO <= x"380030d0"; 
      when 183 => DO <= x"38002061"; 
      when 184 => DO <= x"380030d0"; 
      when 185 => DO <= x"38000000"; 
      when 186 => DO <= x"5f8f892e"; 
      when 187 => DO <= x"4010894b"; 
      when 188 => DO <= x"40108b14"; 
      when 189 => DO <= x"2001905f"; 
      when 190 => DO <= x"4004106f"; 
      when 191 => DO <= x"8bbe200a"; 
      when 192 => DO <= x"001a80ff"; 
      when 193 => DO <= x"60007ff1"; 
      when 194 => DO <= x"84142006"; 
      when 195 => DO <= x"84122005"; 
      when 196 => DO <= x"8b6e2004"; 
      when 197 => DO <= x"8b652006"; 
      when 198 => DO <= x"896e4010"; 
      when 199 => DO <= x"00e48b32"; 
      when 200 => DO <= x"200e8bb5"; 
      when 201 => DO <= x"20028416"; 
      when 202 => DO <= x"2003186f"; 
      when 203 => DO <= x"985f4004"; 
      when 204 => DO <= x"8024200b"; 
      when 205 => DO <= x"044100ea"; 
      when 206 => DO <= x"88bb4010"; 
      when 207 => DO <= x"002105b3"; 
      when 208 => DO <= x"894b4010"; 
      when 209 => DO <= x"89114010"; 
      when 210 => DO <= x"00ba0c3c"; 
      when 211 => DO <= x"00a1508f"; 
      when 212 => DO <= x"30d03800"; 
      when 213 => DO <= x"5e8f10df"; 
      when 214 => DO <= x"905f4014"; 
      when 215 => DO <= x"906f4010"; 
      when 216 => DO <= x"907f400c"; 
      when 217 => DO <= x"908f4008"; 
      when 218 => DO <= x"0c157018"; 
      when 219 => DO <= x"70b1909f"; 
      when 220 => DO <= x"40049085"; 
      when 221 => DO <= x"40089005"; 
      when 222 => DO <= x"40089015"; 
      when 223 => DO <= x"40049815"; 
      when 224 => DO <= x"40048600"; 
      when 225 => DO <= x"60007001"; 
      when 226 => DO <= x"90154024"; 
      when 227 => DO <= x"98154024"; 
      when 228 => DO <= x"90054004"; 
      when 229 => DO <= x"98154004"; 
      when 230 => DO <= x"90054034"; 
      when 231 => DO <= x"98654034"; 
      when 232 => DO <= x"90054014"; 
      when 233 => DO <= x"800e7000"; 
      when 234 => DO <= x"7bb19875"; 
      when 235 => DO <= x"4014c06d"; 
      when 236 => DO <= x"40073800"; 
      when 237 => DO <= x"0c61c36d"; 
      when 238 => DO <= x"40073800"; 
      when 239 => DO <= x"800e7000"; 
      when 240 => DO <= x"7cc1cf2d"; 
      when 241 => DO <= x"40063800"; 
      when 242 => DO <= x"80ff6000"; 
      when 243 => DO <= x"7ff10471"; 
      when 244 => DO <= x"c80d4008"; 
      when 245 => DO <= x"3800800f"; 
      when 246 => DO <= x"70007e91"; 
      when 247 => DO <= x"cd8d4006"; 
      when 248 => DO <= x"38009005"; 
      when 249 => DO <= x"4034800e"; 
      when 250 => DO <= x"70007d51"; 
      when 251 => DO <= x"98754034"; 
      when 252 => DO <= x"cc4d4006"; 
      when 253 => DO <= x"38000c71"; 
      when 254 => DO <= x"cf4d4006"; 
      when 255 => DO <= x"38008afa"; 
      when 256 => DO <= x"60626d57"; 
      when 257 => DO <= x"c0804200"; 
      when 258 => DO <= x"3800ca20"; 
      when 259 => DO <= x"40003800"; 
      when 260 => DO <= x"90054034"; 
      when 261 => DO <= x"800e7000"; 
      when 262 => DO <= x"7f019875"; 
      when 263 => DO <= x"4034c96d"; 
      when 264 => DO <= x"40063800"; 
      when 265 => DO <= x"0c71cc6d"; 
      when 266 => DO <= x"40063800"; 
      when 267 => DO <= x"800f7000"; 
      when 268 => DO <= x"7031c82d"; 
      when 269 => DO <= x"40063800"; 
      when 270 => DO <= x"70096006"; 
      when 271 => DO <= x"c0404200"; 
      when 272 => DO <= x"38007008"; 
      when 273 => DO <= x"cf6d40fc"; 
      when 274 => DO <= x"38006006"; 
      when 275 => DO <= x"c7004200"; 
      when 276 => DO <= x"3800aaaa"; 
      when 277 => DO <= x"70557aa7"; 
      when 278 => DO <= x"0c619005"; 
      when 279 => DO <= x"40345ff1"; 
      when 280 => DO <= x"98254034"; 
      when 281 => DO <= x"10295049"; 
      when 282 => DO <= x"60010627"; 
      when 283 => DO <= x"cea041ff"; 
      when 284 => DO <= x"3800800f"; 
      when 285 => DO <= x"700070e1"; 
      when 286 => DO <= x"c3cd4006"; 
      when 287 => DO <= x"38000c71"; 
      when 288 => DO <= x"c6cd4006"; 
      when 289 => DO <= x"3800aaaa"; 
      when 290 => DO <= x"70557aa7"; 
      when 291 => DO <= x"6006c060"; 
      when 292 => DO <= x"41003800"; 
      when 293 => DO <= x"44c03800"; 
      when 294 => DO <= x"70010c62"; 
      when 295 => DO <= x"18315041"; 
      when 296 => DO <= x"5ff26002"; 
      when 297 => DO <= x"0637cf20"; 
      when 298 => DO <= x"41ff3800"; 
      when 299 => DO <= x"43603800"; 
      when 300 => DO <= x"800e7000"; 
      when 301 => DO <= x"7e31cfed"; 
      when 302 => DO <= x"40053800"; 
      when 303 => DO <= x"4fe03800"; 
      when 304 => DO <= x"800f7000"; 
      when 305 => DO <= x"70e1ceed"; 
      when 306 => DO <= x"40053800"; 
      when 307 => DO <= x"aaaa7055"; 
      when 308 => DO <= x"7aa1aaaa"; 
      when 309 => DO <= x"70557aa7"; 
      when 310 => DO <= x"c14d4006"; 
      when 311 => DO <= x"38004040"; 
      when 312 => DO <= x"38007018"; 
      when 313 => DO <= x"800f7000"; 
      when 314 => DO <= x"71b1ccad"; 
      when 315 => DO <= x"40053800"; 
      when 316 => DO <= x"0c71cfad"; 
      when 317 => DO <= x"40053800"; 
      when 318 => DO <= x"701170b2"; 
      when 319 => DO <= x"90154008"; 
      when 320 => DO <= x"90054008"; 
      when 321 => DO <= x"90254004"; 
      when 322 => DO <= x"04819825"; 
      when 323 => DO <= x"40046001"; 
      when 324 => DO <= x"86006000"; 
      when 325 => DO <= x"70e29025"; 
      when 326 => DO <= x"40249825"; 
      when 327 => DO <= x"40249005"; 
      when 328 => DO <= x"40049825"; 
      when 329 => DO <= x"4004c6a0"; 
      when 330 => DO <= x"41003800"; 
      when 331 => DO <= x"70079005"; 
      when 332 => DO <= x"40349885"; 
      when 333 => DO <= x"40341817"; 
      when 334 => DO <= x"0781c4a0"; 
      when 335 => DO <= x"42003800"; 
      when 336 => DO <= x"800f7000"; 
      when 337 => DO <= x"7241c6ed"; 
      when 338 => DO <= x"40053800"; 
      when 339 => DO <= x"0c71c9ed"; 
      when 340 => DO <= x"40053800"; 
      when 341 => DO <= x"800f7000"; 
      when 342 => DO <= x"73b1c5ad"; 
      when 343 => DO <= x"40053800"; 
      when 344 => DO <= x"0c81c8ad"; 
      when 345 => DO <= x"40053800"; 
      when 346 => DO <= x"800f7000"; 
      when 347 => DO <= x"7481c46d"; 
      when 348 => DO <= x"40053800"; 
      when 349 => DO <= x"1817c76d"; 
      when 350 => DO <= x"40053800"; 
      when 351 => DO <= x"800f7000"; 
      when 352 => DO <= x"7e91c32d"; 
      when 353 => DO <= x"40053800"; 
      when 354 => DO <= x"50475ff6"; 
      when 355 => DO <= x"6006c9c0"; 
      when 356 => DO <= x"41ff3800"; 
      when 357 => DO <= x"800f7000"; 
      when 358 => DO <= x"7501c1ad"; 
      when 359 => DO <= x"40053800"; 
      when 360 => DO <= x"c9ad40fb"; 
      when 361 => DO <= x"3800cb2d"; 
      when 362 => DO <= x"40fb3800"; 
      when 363 => DO <= x"800f7000"; 
      when 364 => DO <= x"7581c02d"; 
      when 365 => DO <= x"40053800"; 
      when 366 => DO <= x"1810c32d"; 
      when 367 => DO <= x"40053800"; 
      when 368 => DO <= x"98104004"; 
      when 369 => DO <= x"c28d4005"; 
      when 370 => DO <= x"3800800f"; 
      when 371 => DO <= x"70007e91"; 
      when 372 => DO <= x"ce4d4004"; 
      when 373 => DO <= x"3800800f"; 
      when 374 => DO <= x"700076f1"; 
      when 375 => DO <= x"cd8d4004"; 
      when 376 => DO <= x"38007001"; 
      when 377 => DO <= x"c80d40fb"; 
      when 378 => DO <= x"3800989f"; 
      when 379 => DO <= x"4004988f"; 
      when 380 => DO <= x"4008987f"; 
      when 381 => DO <= x"400c986f"; 
      when 382 => DO <= x"4010985f"; 
      when 383 => DO <= x"401418df"; 
      when 384 => DO <= x"518f30d0"; 
      when 385 => DO <= x"38000000"; 
      when 386 => DO <= x"5f0f800f"; 
      when 387 => DO <= x"70007871"; 
      when 388 => DO <= x"10df905f"; 
      when 389 => DO <= x"400c906f"; 
      when 390 => DO <= x"4008907f"; 
      when 391 => DO <= x"4004c96d"; 
      when 392 => DO <= x"40043800"; 
      when 393 => DO <= x"ff114000"; 
      when 394 => DO <= x"8000703e"; 
      when 395 => DO <= x"70028000"; 
      when 396 => DO <= x"70409010"; 
      when 397 => DO <= x"40007011"; 
      when 398 => DO <= x"80007040"; 
      when 399 => DO <= x"90004008"; 
      when 400 => DO <= x"80007040"; 
      when 401 => DO <= x"90104008"; 
      when 402 => DO <= x"80007040"; 
      when 403 => DO <= x"90004008"; 
      when 404 => DO <= x"80007040"; 
      when 405 => DO <= x"90204034"; 
      when 406 => DO <= x"80007040"; 
      when 407 => DO <= x"98504034"; 
      when 408 => DO <= x"80007040"; 
      when 409 => DO <= x"90104008"; 
      when 410 => DO <= x"800f7000"; 
      when 411 => DO <= x"7a11c46d"; 
      when 412 => DO <= x"40043800"; 
      when 413 => DO <= x"ffff6001"; 
      when 414 => DO <= x"7ff10451"; 
      when 415 => DO <= x"c70d4004"; 
      when 416 => DO <= x"3800800f"; 
      when 417 => DO <= x"70007e91"; 
      when 418 => DO <= x"c2cd4004"; 
      when 419 => DO <= x"3800800f"; 
      when 420 => DO <= x"70007be1"; 
      when 421 => DO <= x"c20d4004"; 
      when 422 => DO <= x"3800c38d"; 
      when 423 => DO <= x"40fc3800"; 
      when 424 => DO <= x"c4cd4004"; 
      when 425 => DO <= x"3800800f"; 
      when 426 => DO <= x"70007ea1"; 
      when 427 => DO <= x"c08d4004"; 
      when 428 => DO <= x"3800800f"; 
      when 429 => DO <= x"70007ce1"; 
      when 430 => DO <= x"cfcd4003"; 
      when 431 => DO <= x"3800c1cd"; 
      when 432 => DO <= x"40fc3800"; 
      when 433 => DO <= x"c28d4004"; 
      when 434 => DO <= x"3800800f"; 
      when 435 => DO <= x"70007ea1"; 
      when 436 => DO <= x"ce4d4003"; 
      when 437 => DO <= x"3800c96d"; 
      when 438 => DO <= x"40fb3800"; 
      when 439 => DO <= x"0c158956"; 
      when 440 => DO <= x"40106006"; 
      when 441 => DO <= x"c9604200"; 
      when 442 => DO <= x"3800800f"; 
      when 443 => DO <= x"70007dc1"; 
      when 444 => DO <= x"cc4d4003"; 
      when 445 => DO <= x"380080ff"; 
      when 446 => DO <= x"60007ff7"; 
      when 447 => DO <= x"800f7000"; 
      when 448 => DO <= x"7ec1cb2d"; 
      when 449 => DO <= x"40033800"; 
      when 450 => DO <= x"50150475"; 
      when 451 => DO <= x"0c51c6ed"; 
      when 452 => DO <= x"40fb3800"; 
      when 453 => DO <= x"c78d40fb"; 
      when 454 => DO <= x"3800cd2d"; 
      when 455 => DO <= x"40033800"; 
      when 456 => DO <= x"800e7000"; 
      when 457 => DO <= x"7ff1c8ed"; 
      when 458 => DO <= x"40033800"; 
      when 459 => DO <= x"c78d40fb"; 
      when 460 => DO <= x"3800cbad"; 
      when 461 => DO <= x"40033800"; 
      when 462 => DO <= x"800e7000"; 
      when 463 => DO <= x"7ff1c76d"; 
      when 464 => DO <= x"40033800"; 
      when 465 => DO <= x"c50d40fb"; 
      when 466 => DO <= x"3800ca2d"; 
      when 467 => DO <= x"40033800"; 
      when 468 => DO <= x"800e7000"; 
      when 469 => DO <= x"7ff1c5ed"; 
      when 470 => DO <= x"40033800"; 
      when 471 => DO <= x"c40d40fb"; 
      when 472 => DO <= x"3800c8ad"; 
      when 473 => DO <= x"40033800"; 
      when 474 => DO <= x"800f7000"; 
      when 475 => DO <= x"7e91c46d"; 
      when 476 => DO <= x"40033800"; 
      when 477 => DO <= x"5ff66006"; 
      when 478 => DO <= x"c80041ff"; 
      when 479 => DO <= x"38007011"; 
      when 480 => DO <= x"c4cd40fb"; 
      when 481 => DO <= x"38008000"; 
      when 482 => DO <= x"70407001"; 
      when 483 => DO <= x"cc4d40fb"; 
      when 484 => DO <= x"38004fe0"; 
      when 485 => DO <= x"38000000"; 
      when 486 => DO <= x"5fcf7002"; 
      when 487 => DO <= x"81006000"; 
      when 488 => DO <= x"7003aaaa"; 
      when 489 => DO <= x"70557aa4"; 
      when 490 => DO <= x"fffa4000"; 
      when 491 => DO <= x"105f720b"; 
      when 492 => DO <= x"7201881e"; 
      when 493 => DO <= x"4008051e"; 
      when 494 => DO <= x"88e54010"; 
      when 495 => DO <= x"055e8815"; 
      when 496 => DO <= x"4002064e"; 
      when 497 => DO <= x"002510e5"; 
      when 498 => DO <= x"0c1e5ffe"; 
      when 499 => DO <= x"60010ce1"; 
      when 500 => DO <= x"cde041ff"; 
      when 501 => DO <= x"380084ab"; 
      when 502 => DO <= x"2001881e"; 
      when 503 => DO <= x"400805e1"; 
      when 504 => DO <= x"881e4010"; 
      when 505 => DO <= x"05e18614"; 
      when 506 => DO <= x"200e88b1"; 
      when 507 => DO <= x"40028012"; 
      when 508 => DO <= x"20057011"; 
      when 509 => DO <= x"185507e5"; 
      when 510 => DO <= x"c2004100"; 
      when 511 => DO <= x"38000cb1"; 
      when 512 => DO <= x"5ff1600b"; 
      when 513 => DO <= x"0c1bccc0"; 
      when 514 => DO <= x"41ff3800"; 
      when 515 => DO <= x"7001d802"; 
      when 516 => DO <= x"40005ff3"; 
      when 517 => DO <= x"6003c940"; 
      when 518 => DO <= x"41ff3800"; 
      when 519 => DO <= x"185f504f"; 
      when 520 => DO <= x"30d03800"; 
      when 521 => DO <= x"5f8f10df"; 
      when 522 => DO <= x"905f4004"; 
      when 523 => DO <= x"0c15800f"; 
      when 524 => DO <= x"70007f11"; 
      when 525 => DO <= x"c80d4002"; 
      when 526 => DO <= x"38001815"; 
      when 527 => DO <= x"cb0d4002"; 
      when 528 => DO <= x"3800800f"; 
      when 529 => DO <= x"70007e91"; 
      when 530 => DO <= x"c6cd4002"; 
      when 531 => DO <= x"38008010"; 
      when 532 => DO <= x"70007121"; 
      when 533 => DO <= x"c60d4002"; 
      when 534 => DO <= x"38009815"; 
      when 535 => DO <= x"4004c8ed"; 
      when 536 => DO <= x"40023800"; 
      when 537 => DO <= x"80107000"; 
      when 538 => DO <= x"71d1c4ad"; 
      when 539 => DO <= x"40023800"; 
      when 540 => DO <= x"800f7000"; 
      when 541 => DO <= x"7e91c3ed"; 
      when 542 => DO <= x"40023800"; 
      when 543 => DO <= x"80107000"; 
      when 544 => DO <= x"7191c32d"; 
      when 545 => DO <= x"40023800"; 
      when 546 => DO <= x"98154040"; 
      when 547 => DO <= x"c60d4002"; 
      when 548 => DO <= x"38008010"; 
      when 549 => DO <= x"700071d1"; 
      when 550 => DO <= x"c1cd4002"; 
      when 551 => DO <= x"38008010"; 
      when 552 => DO <= x"700071f1"; 
      when 553 => DO <= x"c10d4002"; 
      when 554 => DO <= x"38009815"; 
      when 555 => DO <= x"403cc3ed"; 
      when 556 => DO <= x"40023800"; 
      when 557 => DO <= x"80107000"; 
      when 558 => DO <= x"71d1cfad"; 
      when 559 => DO <= x"40013800"; 
      when 560 => DO <= x"80107000"; 
      when 561 => DO <= x"7251ceed"; 
      when 562 => DO <= x"40013800"; 
      when 563 => DO <= x"98154038"; 
      when 564 => DO <= x"c1cd4002"; 
      when 565 => DO <= x"38008010"; 
      when 566 => DO <= x"700071d1"; 
      when 567 => DO <= x"cd8d4001"; 
      when 568 => DO <= x"38008010"; 
      when 569 => DO <= x"700072b1"; 
      when 570 => DO <= x"cccd4001"; 
      when 571 => DO <= x"38009815"; 
      when 572 => DO <= x"4034cfad"; 
      when 573 => DO <= x"40013800"; 
      when 574 => DO <= x"80107000"; 
      when 575 => DO <= x"71d1cb6d"; 
      when 576 => DO <= x"40013800"; 
      when 577 => DO <= x"800f7000"; 
      when 578 => DO <= x"7e91caad"; 
      when 579 => DO <= x"40013800"; 
      when 580 => DO <= x"80107000"; 
      when 581 => DO <= x"7311c9ed"; 
      when 582 => DO <= x"40013800"; 
      when 583 => DO <= x"98154030"; 
      when 584 => DO <= x"cccd4001"; 
      when 585 => DO <= x"38008010"; 
      when 586 => DO <= x"700071d1"; 
      when 587 => DO <= x"c88d4001"; 
      when 588 => DO <= x"38008010"; 
      when 589 => DO <= x"70007371"; 
      when 590 => DO <= x"c7cd4001"; 
      when 591 => DO <= x"38009815"; 
      when 592 => DO <= x"402ccaad"; 
      when 593 => DO <= x"40013800"; 
      when 594 => DO <= x"80107000"; 
      when 595 => DO <= x"71d1c66d"; 
      when 596 => DO <= x"40013800"; 
      when 597 => DO <= x"80107000"; 
      when 598 => DO <= x"73d1c5ad"; 
      when 599 => DO <= x"40013800"; 
      when 600 => DO <= x"98154028"; 
      when 601 => DO <= x"c88d4001"; 
      when 602 => DO <= x"38008010"; 
      when 603 => DO <= x"700071d1"; 
      when 604 => DO <= x"c44d4001"; 
      when 605 => DO <= x"38008010"; 
      when 606 => DO <= x"70007431"; 
      when 607 => DO <= x"c38d4001"; 
      when 608 => DO <= x"38009815"; 
      when 609 => DO <= x"4024c66d"; 
      when 610 => DO <= x"40013800"; 
      when 611 => DO <= x"80107000"; 
      when 612 => DO <= x"71d1c22d"; 
      when 613 => DO <= x"40013800"; 
      when 614 => DO <= x"800f7000"; 
      when 615 => DO <= x"7e91c16d"; 
      when 616 => DO <= x"40013800"; 
      when 617 => DO <= x"80107000"; 
      when 618 => DO <= x"7491c0ad"; 
      when 619 => DO <= x"40013800"; 
      when 620 => DO <= x"98154020"; 
      when 621 => DO <= x"c38d4001"; 
      when 622 => DO <= x"38008010"; 
      when 623 => DO <= x"700071d1"; 
      when 624 => DO <= x"cf4d4000"; 
      when 625 => DO <= x"38008010"; 
      when 626 => DO <= x"700074f1"; 
      when 627 => DO <= x"ce8d4000"; 
      when 628 => DO <= x"38009815"; 
      when 629 => DO <= x"401cc16d"; 
      when 630 => DO <= x"40013800"; 
      when 631 => DO <= x"80107000"; 
      when 632 => DO <= x"71d1cd2d"; 
      when 633 => DO <= x"40003800"; 
      when 634 => DO <= x"80107000"; 
      when 635 => DO <= x"7551cc6d"; 
      when 636 => DO <= x"40003800"; 
      when 637 => DO <= x"98154018"; 
      when 638 => DO <= x"cf4d4000"; 
      when 639 => DO <= x"38008010"; 
      when 640 => DO <= x"700071d1"; 
      when 641 => DO <= x"cb0d4000"; 
      when 642 => DO <= x"38008010"; 
      when 643 => DO <= x"700075b1"; 
      when 644 => DO <= x"ca4d4000"; 
      when 645 => DO <= x"38009815"; 
      when 646 => DO <= x"4014cd2d"; 
      when 647 => DO <= x"40003800"; 
      when 648 => DO <= x"80107000"; 
      when 649 => DO <= x"71d1c8ed"; 
      when 650 => DO <= x"40003800"; 
      when 651 => DO <= x"800f7000"; 
      when 652 => DO <= x"7e91c82d"; 
      when 653 => DO <= x"40003800"; 
      when 654 => DO <= x"80107000"; 
      when 655 => DO <= x"7611478d"; 
      when 656 => DO <= x"38009815"; 
      when 657 => DO <= x"4010ca6d"; 
      when 658 => DO <= x"40003800"; 
      when 659 => DO <= x"80107000"; 
      when 660 => DO <= x"71d1464d"; 
      when 661 => DO <= x"38008010"; 
      when 662 => DO <= x"70007671"; 
      when 663 => DO <= x"45ad3800"; 
      when 664 => DO <= x"9815400c"; 
      when 665 => DO <= x"c88d4000"; 
      when 666 => DO <= x"38008010"; 
      when 667 => DO <= x"700071d1"; 
      when 668 => DO <= x"446d3800"; 
      when 669 => DO <= x"80107000"; 
      when 670 => DO <= x"76d143cd"; 
      when 671 => DO <= x"38009815"; 
      when 672 => DO <= x"400846cd"; 
      when 673 => DO <= x"38008010"; 
      when 674 => DO <= x"700071d1"; 
      when 675 => DO <= x"42ad3800"; 
      when 676 => DO <= x"800f7000"; 
      when 677 => DO <= x"7e91420d"; 
      when 678 => DO <= x"3800cc6d"; 
      when 679 => DO <= x"40f73800"; 
      when 680 => DO <= x"ff024000"; 
      when 681 => DO <= x"04216201"; 
      when 682 => DO <= x"c0804100"; 
      when 683 => DO <= x"38001815"; 
      when 684 => DO <= x"50211015"; 
      when 685 => DO <= x"4fe03800"; 
      when 686 => DO <= x"5f8f10df"; 
      when 687 => DO <= x"905f4004"; 
      when 688 => DO <= x"0c151a15"; 
      when 689 => DO <= x"6001c180"; 
      when 690 => DO <= x"42003800"; 
      when 691 => DO <= x"3811c50d"; 
      when 692 => DO <= x"40f63800"; 
      when 693 => DO <= x"9a154001"; 
      when 694 => DO <= x"50156001"; 
      when 695 => DO <= x"cec041ff"; 
      when 696 => DO <= x"3800985f"; 
      when 697 => DO <= x"400418df"; 
      when 698 => DO <= x"508f30d0"; 
      when 699 => DO <= x"38000000"; 
      when 700 => DO <= x"5f0f10df"; 
      when 701 => DO <= x"905f400c"; 
      when 702 => DO <= x"0c15906f"; 
      when 703 => DO <= x"40087306"; 
      when 704 => DO <= x"907f4004"; 
      when 705 => DO <= x"ffff703f"; 
      when 706 => DO <= x"6ff58951"; 
      when 707 => DO <= x"401cc060"; 
      when 708 => DO <= x"4a003800"; 
      when 709 => DO <= x"40803800"; 
      when 710 => DO <= x"05614040"; 
      when 711 => DO <= x"38005371"; 
      when 712 => DO <= x"cfed40f5"; 
      when 713 => DO <= x"38008951"; 
      when 714 => DO <= x"401870f7"; 
      when 715 => DO <= x"88524004"; 
      when 716 => DO <= x"ffff703f"; 
      when 717 => DO <= x"6ff20471"; 
      when 718 => DO <= x"c0604a00"; 
      when 719 => DO <= x"38004080"; 
      when 720 => DO <= x"38000561"; 
      when 721 => DO <= x"40403800"; 
      when 722 => DO <= x"5371cd4d"; 
      when 723 => DO <= x"40f53800"; 
      when 724 => DO <= x"89514014"; 
      when 725 => DO <= x"88524008"; 
      when 726 => DO <= x"ffff703f"; 
      when 727 => DO <= x"6ff20471"; 
      when 728 => DO <= x"c0604a00"; 
      when 729 => DO <= x"38004080"; 
      when 730 => DO <= x"38000561"; 
      when 731 => DO <= x"40403800"; 
      when 732 => DO <= x"5371cacd"; 
      when 733 => DO <= x"40f53800"; 
      when 734 => DO <= x"89514010"; 
      when 735 => DO <= x"8852400c"; 
      when 736 => DO <= x"ffff703f"; 
      when 737 => DO <= x"6ff20471"; 
      when 738 => DO <= x"c0604a00"; 
      when 739 => DO <= x"38004080"; 
      when 740 => DO <= x"38000561"; 
      when 741 => DO <= x"40403800"; 
      when 742 => DO <= x"5371c84d"; 
      when 743 => DO <= x"40f53800"; 
      when 744 => DO <= x"8951400c"; 
      when 745 => DO <= x"88524010"; 
      when 746 => DO <= x"ffff703f"; 
      when 747 => DO <= x"6ff20471"; 
      when 748 => DO <= x"c0604a00"; 
      when 749 => DO <= x"38004080"; 
      when 750 => DO <= x"38000561"; 
      when 751 => DO <= x"40403800"; 
      when 752 => DO <= x"5371c5cd"; 
      when 753 => DO <= x"40f53800"; 
      when 754 => DO <= x"89514008"; 
      when 755 => DO <= x"88524014"; 
      when 756 => DO <= x"ffff703f"; 
      when 757 => DO <= x"6ff20471"; 
      when 758 => DO <= x"c0604a00"; 
      when 759 => DO <= x"38004080"; 
      when 760 => DO <= x"38000561"; 
      when 761 => DO <= x"40403800"; 
      when 762 => DO <= x"5371c34d"; 
      when 763 => DO <= x"40f53800"; 
      when 764 => DO <= x"89514004"; 
      when 765 => DO <= x"88524018"; 
      when 766 => DO <= x"ffff703f"; 
      when 767 => DO <= x"6ff20471"; 
      when 768 => DO <= x"c0604a00"; 
      when 769 => DO <= x"38004080"; 
      when 770 => DO <= x"38000561"; 
      when 771 => DO <= x"40403800"; 
      when 772 => DO <= x"5371c0cd"; 
      when 773 => DO <= x"40f53800"; 
      when 774 => DO <= x"84752001"; 
      when 775 => DO <= x"8852401c"; 
      when 776 => DO <= x"ffff703f"; 
      when 777 => DO <= x"6ff2c060"; 
      when 778 => DO <= x"4a003800"; 
      when 779 => DO <= x"40803800"; 
      when 780 => DO <= x"05614040"; 
      when 781 => DO <= x"38005371"; 
      when 782 => DO <= x"ce6d40f4"; 
      when 783 => DO <= x"3800987f"; 
      when 784 => DO <= x"4004986f"; 
      when 785 => DO <= x"4008985f"; 
      when 786 => DO <= x"400c18df"; 
      when 787 => DO <= x"510f30d0"; 
      when 788 => DO <= x"38000000"; 
      when 789 => DO <= x"5f4f10df"; 
      when 790 => DO <= x"905f4008"; 
      when 791 => DO <= x"0c15906f"; 
      when 792 => DO <= x"40047306"; 
      when 793 => DO <= x"809f6000"; 
      when 794 => DO <= x"6ff58951"; 
      when 795 => DO <= x"400cc060"; 
      when 796 => DO <= x"4a003800"; 
      when 797 => DO <= x"40803800"; 
      when 798 => DO <= x"05614040"; 
      when 799 => DO <= x"38005371"; 
      when 800 => DO <= x"c9ed40f4"; 
      when 801 => DO <= x"38008851"; 
      when 802 => DO <= x"400480ff"; 
      when 803 => DO <= x"60007f02"; 
      when 804 => DO <= x"0412809f"; 
      when 805 => DO <= x"60006ff2"; 
      when 806 => DO <= x"8921400c"; 
      when 807 => DO <= x"c0604a00"; 
      when 808 => DO <= x"38004080"; 
      when 809 => DO <= x"38000561"; 
      when 810 => DO <= x"40403800"; 
      when 811 => DO <= x"5371c70d"; 
      when 812 => DO <= x"40f43800"; 
      when 813 => DO <= x"88514008"; 
      when 814 => DO <= x"80ff6000"; 
      when 815 => DO <= x"70020412"; 
      when 816 => DO <= x"809f6000"; 
      when 817 => DO <= x"6ff28921"; 
      when 818 => DO <= x"400cc060"; 
      when 819 => DO <= x"4a003800"; 
      when 820 => DO <= x"40803800"; 
      when 821 => DO <= x"05614040"; 
      when 822 => DO <= x"38005371"; 
      when 823 => DO <= x"c42d40f4"; 
      when 824 => DO <= x"38008851"; 
      when 825 => DO <= x"400c80f0"; 
      when 826 => DO <= x"60007002"; 
      when 827 => DO <= x"0412809f"; 
      when 828 => DO <= x"60006ff2"; 
      when 829 => DO <= x"8921400c"; 
      when 830 => DO <= x"c0604a00"; 
      when 831 => DO <= x"38004080"; 
      when 832 => DO <= x"38000561"; 
      when 833 => DO <= x"40403800"; 
      when 834 => DO <= x"5371c14d"; 
      when 835 => DO <= x"40f43800"; 
      when 836 => DO <= x"986f4004"; 
      when 837 => DO <= x"985f4008"; 
      when 838 => DO <= x"18df50cf"; 
      when 839 => DO <= x"30d03800"; 
      when 840 => DO <= x"5fcf0c14"; 
      when 841 => DO <= x"70017003"; 
      when 842 => DO <= x"10dfcbad"; 
      when 843 => DO <= x"40f53800"; 
      when 844 => DO <= x"18df504f"; 
      when 845 => DO <= x"30d03800"; 
      when 846 => DO <= x"8b212001"; 
      when 847 => DO <= x"89114010"; 
      when 848 => DO <= x"3c023800"; 
      when 849 => DO <= x"88224010"; 
      when 850 => DO <= x"052130d0"; 
      when 851 => DO <= x"38000000"; 
      when 852 => DO <= x"5fcf0c14"; 
      when 853 => DO <= x"70017003"; 
      when 854 => DO <= x"10dfc8ad"; 
      when 855 => DO <= x"40f53800"; 
      when 856 => DO <= x"18df89c2"; 
      when 857 => DO <= x"40108811"; 
      when 858 => DO <= x"40100521"; 
      when 859 => DO <= x"504f30d0"; 
      when 860 => DO <= x"38000000"; 
      when 861 => DO <= x"00000000"; 
      when 862 => DO <= x"00000000"; 
      when 863 => DO <= x"00000000"; 
      when 864 => DO <= x"00000000"; 
      when 865 => DO <= x"00000000"; 
      when 866 => DO <= x"00000000"; 
      when 867 => DO <= x"00000000"; 
      when 868 => DO <= x"00000000"; 
      when 869 => DO <= x"00000000"; 
      when 870 => DO <= x"00000000"; 
      when 871 => DO <= x"00000000"; 
      when 872 => DO <= x"00000000"; 
      when 873 => DO <= x"00000000"; 
      when 874 => DO <= x"00000000"; 
      when 875 => DO <= x"00000000"; 
      when 876 => DO <= x"00000000"; 
      when 877 => DO <= x"00000000"; 
      when 878 => DO <= x"00000000"; 
      when 879 => DO <= x"00000000"; 
      when 880 => DO <= x"00000000"; 
      when 881 => DO <= x"00000000"; 
      when 882 => DO <= x"00000000"; 
      when 883 => DO <= x"00000000"; 
      when 884 => DO <= x"00000000"; 
      when 885 => DO <= x"00000000"; 
      when 886 => DO <= x"00000000"; 
      when 887 => DO <= x"00000000"; 
      when 888 => DO <= x"00000000"; 
      when 889 => DO <= x"00000000"; 
      when 890 => DO <= x"00000000"; 
      when 891 => DO <= x"00000000"; 
      when 892 => DO <= x"00000000"; 
      when 893 => DO <= x"00000000"; 
      when 894 => DO <= x"00000000"; 
      when 895 => DO <= x"00000000"; 
      when 896 => DO <= x"c88040f3"; 
      when 897 => DO <= x"38000000"; 
      when 898 => DO <= x"00000000"; 
      when 899 => DO <= x"00000000"; 
      when 900 => DO <= x"c78040f3"; 
      when 901 => DO <= x"38000000"; 
      when 902 => DO <= x"00000000"; 
      when 903 => DO <= x"00000000"; 
      when 904 => DO <= x"c68040f3"; 
      when 905 => DO <= x"38000000"; 
      when 906 => DO <= x"00000000"; 
      when 907 => DO <= x"00000000"; 
      when 908 => DO <= x"c58040f3"; 
      when 909 => DO <= x"38000000"; 
      when 910 => DO <= x"00000000"; 
      when 911 => DO <= x"00000000"; 
      when 912 => DO <= x"c48040f3"; 
      when 913 => DO <= x"38000000"; 
      when 914 => DO <= x"4d656d6f"; 
      when 915 => DO <= x"72792065"; 
      when 916 => DO <= x"72726f72"; 
      when 917 => DO <= x"20617420"; 
      when 918 => DO <= x"61646472"; 
      when 919 => DO <= x"65737320"; 
      when 920 => DO <= x"00200058"; 
      when 921 => DO <= x"5468756e"; 
      when 922 => DO <= x"64657243"; 
      when 923 => DO <= x"6f726520"; 
      when 924 => DO <= x"426f6f74"; 
      when 925 => DO <= x"204c6f61"; 
      when 926 => DO <= x"64657220"; 
      when 927 => DO <= x"76302e31"; 
      when 928 => DO <= x"20284329"; 
      when 929 => DO <= x"20323031"; 
      when 930 => DO <= x"3420416c"; 
      when 931 => DO <= x"7661726f"; 
      when 932 => DO <= x"204c6f70"; 
      when 933 => DO <= x"65730d0a"; 
      when 934 => DO <= x"54657374"; 
      when 935 => DO <= x"696e6720"; 
      when 936 => DO <= x"6d656d6f"; 
      when 937 => DO <= x"72793a20"; 
      when 938 => DO <= x"00466169"; 
      when 939 => DO <= x"6c65640d"; 
      when 940 => DO <= x"0a005061"; 
      when 941 => DO <= x"73736564"; 
      when 942 => DO <= x"0d0a0050"; 
      when 943 => DO <= x"726f6772"; 
      when 944 => DO <= x"616d2073"; 
      when 945 => DO <= x"697a653a"; 
      when 946 => DO <= x"20307800"; 
      when 947 => DO <= x"2c204352"; 
      when 948 => DO <= x"43203078"; 
      when 949 => DO <= x"00536967"; 
      when 950 => DO <= x"6e617475"; 
      when 951 => DO <= x"72653a20"; 
      when 952 => DO <= x"30780020"; 
      when 953 => DO <= x"2d20494e"; 
      when 954 => DO <= x"56414c49"; 
      when 955 => DO <= x"440d0a00"; 
      when 956 => DO <= x"0d0a5461"; 
      when 957 => DO <= x"72676574"; 
      when 958 => DO <= x"20626f61"; 
      when 959 => DO <= x"72643a20"; 
      when 960 => DO <= x"3078000d"; 
      when 961 => DO <= x"0a4c6f61"; 
      when 962 => DO <= x"64696e67"; 
      when 963 => DO <= x"3a004368"; 
      when 964 => DO <= x"65636b73"; 
      when 965 => DO <= x"756d3a20"; 
      when 966 => DO <= x"3078002c"; 
      when 967 => DO <= x"206d656d"; 
      when 968 => DO <= x"20307800"; 
      when 969 => DO <= x"4d69736d"; 
      when 970 => DO <= x"61746368"; 
      when 971 => DO <= x"20617420"; 
      when 972 => DO <= x"61646472"; 
      when 973 => DO <= x"65737320"; 
      when 974 => DO <= x"3078002c"; 
      when 975 => DO <= x"20657870"; 
      when 976 => DO <= x"65637469"; 
      when 977 => DO <= x"6e672000"; 
      when 978 => DO <= x"2c207265"; 
      when 979 => DO <= x"61642000"; 
      when 980 => DO <= x"20646f6e"; 
      when 981 => DO <= x"650d0a00"; 
      when 982 => DO <= x"496e6974"; 
      when 983 => DO <= x"69616c20"; 
      when 984 => DO <= x"6d656d6f"; 
      when 985 => DO <= x"72792062"; 
      when 986 => DO <= x"79746573"; 
      when 987 => DO <= x"3a200053"; 
      when 988 => DO <= x"74617274"; 
      when 989 => DO <= x"696e6720"; 
      when 990 => DO <= x"6170706c"; 
      when 991 => DO <= x"69636174"; 
      when 992 => DO <= x"696f6e2e"; 
      when 993 => DO <= x"0d0a0043"; 
      when 994 => DO <= x"6f6e6e65"; 
      when 995 => DO <= x"6374696e"; 
      when 996 => DO <= x"6720746f"; 
      when 997 => DO <= x"20535049"; 
      when 998 => DO <= x"20666c61"; 
      when 999 => DO <= x"73680d0a"; 
      when 1000 => DO <= x"00535049"; 
      when 1001 => DO <= x"20466c61"; 
      when 1002 => DO <= x"73682049"; 
      when 1003 => DO <= x"64656e74"; 
      when 1004 => DO <= x"69666963"; 
      when 1005 => DO <= x"6174696f"; 
      when 1006 => DO <= x"6e3a2030"; 
      when 1007 => DO <= x"78004661"; 
      when 1008 => DO <= x"756c7420"; 
      when 1009 => DO <= x"61646472"; 
      when 1010 => DO <= x"6573733a"; 
      when 1011 => DO <= x"20004661"; 
      when 1012 => DO <= x"756c7420"; 
      when 1013 => DO <= x"666c6167"; 
      when 1014 => DO <= x"733a2000"; 
      when 1015 => DO <= x"54726163"; 
      when 1016 => DO <= x"65627566"; 
      when 1017 => DO <= x"6665723a"; 
      when 1018 => DO <= x"200d0a00"; 
      when 1019 => DO <= x"45203078"; 
      when 1020 => DO <= x"000d0a45"; 
      when 1021 => DO <= x"78636570"; 
      when 1022 => DO <= x"74696f6e"; 
      when 1023 => DO <= x"20636175"; 
      when 1024 => DO <= x"67687420"; 
      when 1025 => DO <= x"61742061"; 
      when 1026 => DO <= x"64647265"; 
      when 1027 => DO <= x"73732030"; 
      when 1028 => DO <= x"78005350"; 
      when 1029 => DO <= x"53523a20"; 
      when 1030 => DO <= x"00523120"; 
      when 1031 => DO <= x"3a200052"; 
      when 1032 => DO <= x"32203a20"; 
      when 1033 => DO <= x"00523320"; 
      when 1034 => DO <= x"3a200052"; 
      when 1035 => DO <= x"34203a20"; 
      when 1036 => DO <= x"00523520"; 
      when 1037 => DO <= x"3a200052"; 
      when 1038 => DO <= x"36203a20"; 
      when 1039 => DO <= x"00523720"; 
      when 1040 => DO <= x"3a200052"; 
      when 1041 => DO <= x"38203a20"; 
      when 1042 => DO <= x"00523920"; 
      when 1043 => DO <= x"3a200052"; 
      when 1044 => DO <= x"31303a20"; 
      when 1045 => DO <= x"00523131"; 
      when 1046 => DO <= x"3a200052"; 
      when 1047 => DO <= x"31323a20"; 
      when 1048 => DO <= x"00523133"; 
      when 1049 => DO <= x"3a200052"; 
      when 1050 => DO <= x"31343a20"; 
      when 1051 => DO <= x"00523135"; 
      when 1052 => DO <= x"3a200000"; 
      when 1053 => DO <= x"00000000"; 
      when 1054 => DO <= x"12345678"; 
      when 1055 => DO <= x"00000002"; 
      when 1056 => DO <= x"00000000"; 
      when 1057 => DO <= x"00000000"; 
      when 1058 => DO <= x"00000000"; 
      when 1059 => DO <= x"00000000"; 
      when 1060 => DO <= x"00000000"; 
      when 1061 => DO <= x"00000000"; 
      when 1062 => DO <= x"00000000"; 
      when 1063 => DO <= x"00000000"; 
      when 1064 => DO <= x"00000000"; 
      when 1065 => DO <= x"00000000"; 
      when 1066 => DO <= x"00000000"; 
      when 1067 => DO <= x"00000000"; 
      when 1068 => DO <= x"00000000"; 
      when 1069 => DO <= x"00000000"; 
      when 1070 => DO <= x"00000000"; 
      when 1071 => DO <= x"00000000"; 
      when 1072 => DO <= x"00000000"; 
      when 1073 => DO <= x"00000000"; 
      when 1074 => DO <= x"00000000"; 
      when 1075 => DO <= x"00000000"; 
      when 1076 => DO <= x"00000000"; 
      when 1077 => DO <= x"00000000"; 
      when 1078 => DO <= x"00000000"; 
      when 1079 => DO <= x"00000000"; 
      when 1080 => DO <= x"00000000"; 
      when 1081 => DO <= x"00000000"; 
      when 1082 => DO <= x"00000000"; 
      when 1083 => DO <= x"00000000"; 
      when 1084 => DO <= x"00000000"; 
      when 1085 => DO <= x"00000000"; 
      when 1086 => DO <= x"00000000"; 
      when 1087 => DO <= x"00000000"; 
      when 1088 => DO <= x"00000000"; 
      when 1089 => DO <= x"00000000"; 
      when 1090 => DO <= x"00000000"; 
      when 1091 => DO <= x"00000000"; 
      when 1092 => DO <= x"00000000"; 
      when 1093 => DO <= x"00000000"; 
      when 1094 => DO <= x"00000000"; 
      when 1095 => DO <= x"00000000"; 
      when 1096 => DO <= x"00000000"; 
      when 1097 => DO <= x"00000000"; 
      when 1098 => DO <= x"00000000"; 
      when 1099 => DO <= x"00000000"; 
      when 1100 => DO <= x"00000000"; 
      when 1101 => DO <= x"00000000"; 
      when 1102 => DO <= x"00000000"; 
      when 1103 => DO <= x"00000000"; 
      when 1104 => DO <= x"00000000"; 
      when 1105 => DO <= x"00000000"; 
      when 1106 => DO <= x"00000000"; 
      when 1107 => DO <= x"00000000"; 
      when 1108 => DO <= x"00000000"; 
      when 1109 => DO <= x"00000000"; 
      when 1110 => DO <= x"00000000"; 
      when 1111 => DO <= x"00000000"; 
      when 1112 => DO <= x"00000000"; 
      when 1113 => DO <= x"00000000"; 
      when 1114 => DO <= x"00000000"; 
      when 1115 => DO <= x"00000000"; 
      when 1116 => DO <= x"00000000"; 
      when 1117 => DO <= x"00000000"; 
      when 1118 => DO <= x"00000000"; 
      when 1119 => DO <= x"00000000"; 
      when 1120 => DO <= x"00000000"; 
      when 1121 => DO <= x"00000000"; 
      when 1122 => DO <= x"00000000"; 
      when 1123 => DO <= x"00000000"; 
      when 1124 => DO <= x"00000000"; 
      when 1125 => DO <= x"00000000"; 
      when 1126 => DO <= x"00000000"; 
      when 1127 => DO <= x"00000000"; 
      when 1128 => DO <= x"00000000"; 
      when 1129 => DO <= x"00000000"; 
      when 1130 => DO <= x"00000000"; 
      when 1131 => DO <= x"00000000"; 
      when 1132 => DO <= x"00000000"; 
      when 1133 => DO <= x"00000000"; 
      when 1134 => DO <= x"00000000"; 
      when 1135 => DO <= x"00000000"; 
      when 1136 => DO <= x"00000000"; 
      when 1137 => DO <= x"00000000"; 
      when 1138 => DO <= x"00000000"; 
      when 1139 => DO <= x"00000000"; 
      when 1140 => DO <= x"00000000"; 
      when 1141 => DO <= x"00000000"; 
      when 1142 => DO <= x"00000000"; 
      when 1143 => DO <= x"00000000"; 
      when 1144 => DO <= x"00000000"; 
      when 1145 => DO <= x"00000000"; 
      when 1146 => DO <= x"00000000"; 
      when 1147 => DO <= x"00000000"; 
      when 1148 => DO <= x"00000000"; 
      when 1149 => DO <= x"00000000"; 
      when 1150 => DO <= x"00000000"; 
      when 1151 => DO <= x"00000000"; 
      when 1152 => DO <= x"00000000"; 
      when 1153 => DO <= x"00000000"; 
      when 1154 => DO <= x"00000000"; 
      when 1155 => DO <= x"00000000"; 
      when 1156 => DO <= x"00000000"; 
      when 1157 => DO <= x"00000000"; 
      when 1158 => DO <= x"00000000"; 
      when 1159 => DO <= x"00000000"; 
      when 1160 => DO <= x"00000000"; 
      when 1161 => DO <= x"00000000"; 
      when 1162 => DO <= x"00000000"; 
      when 1163 => DO <= x"00000000"; 
      when 1164 => DO <= x"00000000"; 
      when 1165 => DO <= x"00000000"; 
      when 1166 => DO <= x"00000000"; 
      when 1167 => DO <= x"00000000"; 
      when 1168 => DO <= x"00000000"; 
      when 1169 => DO <= x"00000000"; 
      when 1170 => DO <= x"00000000"; 
      when 1171 => DO <= x"00000000"; 
      when 1172 => DO <= x"00000000"; 
      when 1173 => DO <= x"00000000"; 
      when 1174 => DO <= x"00000000"; 
      when 1175 => DO <= x"00000000"; 
      when 1176 => DO <= x"00000000"; 
      when 1177 => DO <= x"00000000"; 
      when 1178 => DO <= x"00000000"; 
      when 1179 => DO <= x"00000000"; 
      when 1180 => DO <= x"00000000"; 
      when 1181 => DO <= x"00000000"; 
      when 1182 => DO <= x"00000000"; 
      when 1183 => DO <= x"00000000"; 
      when 1184 => DO <= x"00000000"; 
      when 1185 => DO <= x"00000000"; 
      when 1186 => DO <= x"00000000"; 
      when 1187 => DO <= x"00000000"; 
      when 1188 => DO <= x"00000000"; 
      when 1189 => DO <= x"00000000"; 
      when 1190 => DO <= x"00000000"; 
      when 1191 => DO <= x"00000000"; 
      when 1192 => DO <= x"00000000"; 
      when 1193 => DO <= x"00000000"; 
      when 1194 => DO <= x"00000000"; 
      when 1195 => DO <= x"00000000"; 
      when 1196 => DO <= x"00000000"; 
      when 1197 => DO <= x"00000000"; 
      when 1198 => DO <= x"00000000"; 
      when 1199 => DO <= x"00000000"; 
      when 1200 => DO <= x"00000000"; 
      when 1201 => DO <= x"00000000"; 
      when 1202 => DO <= x"00000000"; 
      when 1203 => DO <= x"00000000"; 
      when 1204 => DO <= x"00000000"; 
      when 1205 => DO <= x"00000000"; 
      when 1206 => DO <= x"00000000"; 
      when 1207 => DO <= x"00000000"; 
      when 1208 => DO <= x"00000000"; 
      when 1209 => DO <= x"00000000"; 
      when 1210 => DO <= x"00000000"; 
      when 1211 => DO <= x"00000000"; 
      when 1212 => DO <= x"00000000"; 
      when 1213 => DO <= x"00000000"; 
      when 1214 => DO <= x"00000000"; 
      when 1215 => DO <= x"00000000"; 
      when 1216 => DO <= x"00000000"; 
      when 1217 => DO <= x"00000000"; 
      when 1218 => DO <= x"00000000"; 
      when 1219 => DO <= x"00000000"; 
      when 1220 => DO <= x"00000000"; 
      when 1221 => DO <= x"00000000"; 
      when 1222 => DO <= x"00000000"; 
      when 1223 => DO <= x"00000000"; 
      when 1224 => DO <= x"00000000"; 
      when 1225 => DO <= x"00000000"; 
      when 1226 => DO <= x"00000000"; 
      when 1227 => DO <= x"00000000"; 
      when 1228 => DO <= x"00000000"; 
      when 1229 => DO <= x"00000000"; 
      when 1230 => DO <= x"00000000"; 
      when 1231 => DO <= x"00000000"; 
      when 1232 => DO <= x"00000000"; 
      when 1233 => DO <= x"00000000"; 
      when 1234 => DO <= x"00000000"; 
      when 1235 => DO <= x"00000000"; 
      when 1236 => DO <= x"00000000"; 
      when 1237 => DO <= x"00000000"; 
      when 1238 => DO <= x"00000000"; 
      when 1239 => DO <= x"00000000"; 
      when 1240 => DO <= x"00000000"; 
      when 1241 => DO <= x"00000000"; 
      when 1242 => DO <= x"00000000"; 
      when 1243 => DO <= x"00000000"; 
      when 1244 => DO <= x"00000000"; 
      when 1245 => DO <= x"00000000"; 
      when 1246 => DO <= x"00000000"; 
      when 1247 => DO <= x"00000000"; 
      when 1248 => DO <= x"00000000"; 
      when 1249 => DO <= x"00000000"; 
      when 1250 => DO <= x"00000000"; 
      when 1251 => DO <= x"00000000"; 
      when 1252 => DO <= x"00000000"; 
      when 1253 => DO <= x"00000000"; 
      when 1254 => DO <= x"00000000"; 
      when 1255 => DO <= x"00000000"; 
      when 1256 => DO <= x"00000000"; 
      when 1257 => DO <= x"00000000"; 
      when 1258 => DO <= x"00000000"; 
      when 1259 => DO <= x"00000000"; 
      when 1260 => DO <= x"00000000"; 
      when 1261 => DO <= x"00000000"; 
      when 1262 => DO <= x"00000000"; 
      when 1263 => DO <= x"00000000"; 
      when 1264 => DO <= x"00000000"; 
      when 1265 => DO <= x"00000000"; 
      when 1266 => DO <= x"00000000"; 
      when 1267 => DO <= x"00000000"; 
      when 1268 => DO <= x"00000000"; 
      when 1269 => DO <= x"00000000"; 
      when 1270 => DO <= x"00000000"; 
      when 1271 => DO <= x"00000000"; 
      when 1272 => DO <= x"00000000"; 
      when 1273 => DO <= x"00000000"; 
      when 1274 => DO <= x"00000000"; 
      when 1275 => DO <= x"00000000"; 
      when 1276 => DO <= x"00000000"; 
      when 1277 => DO <= x"00000000"; 
      when 1278 => DO <= x"00000000"; 
      when 1279 => DO <= x"00000000"; 
      when 1280 => DO <= x"00000000"; 
      when 1281 => DO <= x"00000000"; 
      when 1282 => DO <= x"00000000"; 
      when 1283 => DO <= x"00000000"; 
      when 1284 => DO <= x"00000000"; 
      when 1285 => DO <= x"00000000"; 
      when 1286 => DO <= x"00000000"; 
      when 1287 => DO <= x"00000000"; 
      when 1288 => DO <= x"00000000"; 
      when 1289 => DO <= x"00000000"; 
      when 1290 => DO <= x"00000000"; 
      when 1291 => DO <= x"00000000"; 
      when 1292 => DO <= x"00000000"; 
      when 1293 => DO <= x"00000000"; 
      when 1294 => DO <= x"00000000"; 
      when 1295 => DO <= x"00000000"; 
      when 1296 => DO <= x"00000000"; 
      when 1297 => DO <= x"00000000"; 
      when 1298 => DO <= x"00000000"; 
      when 1299 => DO <= x"00000000"; 
      when 1300 => DO <= x"00000000"; 
      when 1301 => DO <= x"00000000"; 
      when 1302 => DO <= x"00000000"; 
      when 1303 => DO <= x"00000000"; 
      when 1304 => DO <= x"00000000"; 
      when 1305 => DO <= x"00000000"; 
      when 1306 => DO <= x"00000000"; 
      when 1307 => DO <= x"00000000"; 
      when 1308 => DO <= x"00000000"; 
      when 1309 => DO <= x"00000000"; 
      when 1310 => DO <= x"00000000"; 
      when 1311 => DO <= x"00000000"; 
      when 1312 => DO <= x"00000000"; 
      when 1313 => DO <= x"00000000"; 
      when 1314 => DO <= x"00000000"; 
      when 1315 => DO <= x"00000000"; 
      when 1316 => DO <= x"00000000"; 
      when 1317 => DO <= x"00000000"; 
      when 1318 => DO <= x"00000000"; 
      when 1319 => DO <= x"00000000"; 
      when 1320 => DO <= x"00000000"; 
      when 1321 => DO <= x"00000000"; 
      when 1322 => DO <= x"00000000"; 
      when 1323 => DO <= x"00000000"; 
      when 1324 => DO <= x"00000000"; 
      when 1325 => DO <= x"00000000"; 
      when 1326 => DO <= x"00000000"; 
      when 1327 => DO <= x"00000000"; 
      when 1328 => DO <= x"00000000"; 
      when 1329 => DO <= x"00000000"; 
      when 1330 => DO <= x"00000000"; 
      when 1331 => DO <= x"00000000"; 
      when 1332 => DO <= x"00000000"; 
      when 1333 => DO <= x"00000000"; 
      when 1334 => DO <= x"00000000"; 
      when 1335 => DO <= x"00000000"; 
      when 1336 => DO <= x"00000000"; 
      when 1337 => DO <= x"00000000"; 
      when 1338 => DO <= x"00000000"; 
      when 1339 => DO <= x"00000000"; 
      when 1340 => DO <= x"00000000"; 
      when 1341 => DO <= x"00000000"; 
      when 1342 => DO <= x"00000000"; 
      when 1343 => DO <= x"00000000"; 
      when 1344 => DO <= x"00000000"; 
      when 1345 => DO <= x"00000000"; 
      when 1346 => DO <= x"00000000"; 
      when 1347 => DO <= x"00000000"; 
      when 1348 => DO <= x"00000000"; 
      when 1349 => DO <= x"00000000"; 
      when 1350 => DO <= x"00000000"; 
      when 1351 => DO <= x"00000000"; 
      when 1352 => DO <= x"00000000"; 
      when 1353 => DO <= x"00000000"; 
      when 1354 => DO <= x"00000000"; 
      when 1355 => DO <= x"00000000"; 
      when 1356 => DO <= x"00000000"; 
      when 1357 => DO <= x"00000000"; 
      when 1358 => DO <= x"00000000"; 
      when 1359 => DO <= x"00000000"; 
      when 1360 => DO <= x"00000000"; 
      when 1361 => DO <= x"00000000"; 
      when 1362 => DO <= x"00000000"; 
      when 1363 => DO <= x"00000000"; 
      when 1364 => DO <= x"00000000"; 
      when 1365 => DO <= x"00000000"; 
      when 1366 => DO <= x"00000000"; 
      when 1367 => DO <= x"00000000"; 
      when 1368 => DO <= x"00000000"; 
      when 1369 => DO <= x"00000000"; 
      when 1370 => DO <= x"00000000"; 
      when 1371 => DO <= x"00000000"; 
      when 1372 => DO <= x"00000000"; 
      when 1373 => DO <= x"00000000"; 
      when 1374 => DO <= x"00000000"; 
      when 1375 => DO <= x"00000000"; 
      when 1376 => DO <= x"00000000"; 
      when 1377 => DO <= x"00000000"; 
      when 1378 => DO <= x"00000000"; 
      when 1379 => DO <= x"00000000"; 
      when 1380 => DO <= x"00000000"; 
      when 1381 => DO <= x"00000000"; 
      when 1382 => DO <= x"00000000"; 
      when 1383 => DO <= x"00000000"; 
      when 1384 => DO <= x"00000000"; 
      when 1385 => DO <= x"00000000"; 
      when 1386 => DO <= x"00000000"; 
      when 1387 => DO <= x"00000000"; 
      when 1388 => DO <= x"00000000"; 
      when 1389 => DO <= x"00000000"; 
      when 1390 => DO <= x"00000000"; 
      when 1391 => DO <= x"00000000"; 
      when 1392 => DO <= x"00000000"; 
      when 1393 => DO <= x"00000000"; 
      when 1394 => DO <= x"00000000"; 
      when 1395 => DO <= x"00000000"; 
      when 1396 => DO <= x"00000000"; 
      when 1397 => DO <= x"00000000"; 
      when 1398 => DO <= x"00000000"; 
      when 1399 => DO <= x"00000000"; 
      when 1400 => DO <= x"00000000"; 
      when 1401 => DO <= x"00000000"; 
      when 1402 => DO <= x"00000000"; 
      when 1403 => DO <= x"00000000"; 
      when 1404 => DO <= x"00000000"; 
      when 1405 => DO <= x"00000000"; 
      when 1406 => DO <= x"00000000"; 
      when 1407 => DO <= x"00000000"; 
      when 1408 => DO <= x"00000000"; 
      when 1409 => DO <= x"00000000"; 
      when 1410 => DO <= x"00000000"; 
      when 1411 => DO <= x"00000000"; 
      when 1412 => DO <= x"00000000"; 
      when 1413 => DO <= x"00000000"; 
      when 1414 => DO <= x"00000000"; 
      when 1415 => DO <= x"00000000"; 
      when 1416 => DO <= x"00000000"; 
      when 1417 => DO <= x"00000000"; 
      when 1418 => DO <= x"00000000"; 
      when 1419 => DO <= x"00000000"; 
      when 1420 => DO <= x"00000000"; 
      when 1421 => DO <= x"00000000"; 
      when 1422 => DO <= x"00000000"; 
      when 1423 => DO <= x"00000000"; 
      when 1424 => DO <= x"00000000"; 
      when 1425 => DO <= x"00000000"; 
      when 1426 => DO <= x"00000000"; 
      when 1427 => DO <= x"00000000"; 
      when 1428 => DO <= x"00000000"; 
      when 1429 => DO <= x"00000000"; 
      when 1430 => DO <= x"00000000"; 
      when 1431 => DO <= x"00000000"; 
      when 1432 => DO <= x"00000000"; 
      when 1433 => DO <= x"00000000"; 
      when 1434 => DO <= x"00000000"; 
      when 1435 => DO <= x"00000000"; 
      when 1436 => DO <= x"00000000"; 
      when 1437 => DO <= x"00000000"; 
      when 1438 => DO <= x"00000000"; 
      when 1439 => DO <= x"00000000"; 
      when 1440 => DO <= x"00000000"; 
      when 1441 => DO <= x"00000000"; 
      when 1442 => DO <= x"00000000"; 
      when 1443 => DO <= x"00000000"; 
      when 1444 => DO <= x"00000000"; 
      when 1445 => DO <= x"00000000"; 
      when 1446 => DO <= x"00000000"; 
      when 1447 => DO <= x"00000000"; 
      when 1448 => DO <= x"00000000"; 
      when 1449 => DO <= x"00000000"; 
      when 1450 => DO <= x"00000000"; 
      when 1451 => DO <= x"00000000"; 
      when 1452 => DO <= x"00000000"; 
      when 1453 => DO <= x"00000000"; 
      when 1454 => DO <= x"00000000"; 
      when 1455 => DO <= x"00000000"; 
      when 1456 => DO <= x"00000000"; 
      when 1457 => DO <= x"00000000"; 
      when 1458 => DO <= x"00000000"; 
      when 1459 => DO <= x"00000000"; 
      when 1460 => DO <= x"00000000"; 
      when 1461 => DO <= x"00000000"; 
      when 1462 => DO <= x"00000000"; 
      when 1463 => DO <= x"00000000"; 
      when 1464 => DO <= x"00000000"; 
      when 1465 => DO <= x"00000000"; 
      when 1466 => DO <= x"00000000"; 
      when 1467 => DO <= x"00000000"; 
      when 1468 => DO <= x"00000000"; 
      when 1469 => DO <= x"00000000"; 
      when 1470 => DO <= x"00000000"; 
      when 1471 => DO <= x"00000000"; 
      when 1472 => DO <= x"00000000"; 
      when 1473 => DO <= x"00000000"; 
      when 1474 => DO <= x"00000000"; 
      when 1475 => DO <= x"00000000"; 
      when 1476 => DO <= x"00000000"; 
      when 1477 => DO <= x"00000000"; 
      when 1478 => DO <= x"00000000"; 
      when 1479 => DO <= x"00000000"; 
      when 1480 => DO <= x"00000000"; 
      when 1481 => DO <= x"00000000"; 
      when 1482 => DO <= x"00000000"; 
      when 1483 => DO <= x"00000000"; 
      when 1484 => DO <= x"00000000"; 
      when 1485 => DO <= x"00000000"; 
      when 1486 => DO <= x"00000000"; 
      when 1487 => DO <= x"00000000"; 
      when 1488 => DO <= x"00000000"; 
      when 1489 => DO <= x"00000000"; 
      when 1490 => DO <= x"00000000"; 
      when 1491 => DO <= x"00000000"; 
      when 1492 => DO <= x"00000000"; 
      when 1493 => DO <= x"00000000"; 
      when 1494 => DO <= x"00000000"; 
      when 1495 => DO <= x"00000000"; 
      when 1496 => DO <= x"00000000"; 
      when 1497 => DO <= x"00000000"; 
      when 1498 => DO <= x"00000000"; 
      when 1499 => DO <= x"00000000"; 
      when 1500 => DO <= x"00000000"; 
      when 1501 => DO <= x"00000000"; 
      when 1502 => DO <= x"00000000"; 
      when 1503 => DO <= x"00000000"; 
      when 1504 => DO <= x"00000000"; 
      when 1505 => DO <= x"00000000"; 
      when 1506 => DO <= x"00000000"; 
      when 1507 => DO <= x"00000000"; 
      when 1508 => DO <= x"00000000"; 
      when 1509 => DO <= x"00000000"; 
      when 1510 => DO <= x"00000000"; 
      when 1511 => DO <= x"00000000"; 
      when 1512 => DO <= x"00000000"; 
      when 1513 => DO <= x"00000000"; 
      when 1514 => DO <= x"00000000"; 
      when 1515 => DO <= x"00000000"; 
      when 1516 => DO <= x"00000000"; 
      when 1517 => DO <= x"00000000"; 
      when 1518 => DO <= x"00000000"; 
      when 1519 => DO <= x"00000000"; 
      when 1520 => DO <= x"00000000"; 
      when 1521 => DO <= x"00000000"; 
      when 1522 => DO <= x"00000000"; 
      when 1523 => DO <= x"00000000"; 
      when 1524 => DO <= x"00000000"; 
      when 1525 => DO <= x"00000000"; 
      when 1526 => DO <= x"00000000"; 
      when 1527 => DO <= x"00000000"; 
      when 1528 => DO <= x"00000000"; 
      when 1529 => DO <= x"00000000"; 
      when 1530 => DO <= x"00000000"; 
      when 1531 => DO <= x"00000000"; 
      when 1532 => DO <= x"00000000"; 
      when 1533 => DO <= x"00000000"; 
      when 1534 => DO <= x"00000000"; 
      when 1535 => DO <= x"00000000"; 
      when 1536 => DO <= x"00000000"; 
      when 1537 => DO <= x"00000000"; 
      when 1538 => DO <= x"00000000"; 
      when 1539 => DO <= x"00000000"; 
      when 1540 => DO <= x"00000000"; 
      when 1541 => DO <= x"00000000"; 
      when 1542 => DO <= x"00000000"; 
      when 1543 => DO <= x"00000000"; 
      when 1544 => DO <= x"00000000"; 
      when 1545 => DO <= x"00000000"; 
      when 1546 => DO <= x"00000000"; 
      when 1547 => DO <= x"00000000"; 
      when 1548 => DO <= x"00000000"; 
      when 1549 => DO <= x"00000000"; 
      when 1550 => DO <= x"00000000"; 
      when 1551 => DO <= x"00000000"; 
      when 1552 => DO <= x"00000000"; 
      when 1553 => DO <= x"00000000"; 
      when 1554 => DO <= x"00000000"; 
      when 1555 => DO <= x"00000000"; 
      when 1556 => DO <= x"00000000"; 
      when 1557 => DO <= x"00000000"; 
      when 1558 => DO <= x"00000000"; 
      when 1559 => DO <= x"00000000"; 
      when 1560 => DO <= x"00000000"; 
      when 1561 => DO <= x"00000000"; 
      when 1562 => DO <= x"00000000"; 
      when 1563 => DO <= x"00000000"; 
      when 1564 => DO <= x"00000000"; 
      when 1565 => DO <= x"00000000"; 
      when 1566 => DO <= x"00000000"; 
      when 1567 => DO <= x"00000000"; 
      when 1568 => DO <= x"00000000"; 
      when 1569 => DO <= x"00000000"; 
      when 1570 => DO <= x"00000000"; 
      when 1571 => DO <= x"00000000"; 
      when 1572 => DO <= x"00000000"; 
      when 1573 => DO <= x"00000000"; 
      when 1574 => DO <= x"00000000"; 
      when 1575 => DO <= x"00000000"; 
      when 1576 => DO <= x"00000000"; 
      when 1577 => DO <= x"00000000"; 
      when 1578 => DO <= x"00000000"; 
      when 1579 => DO <= x"00000000"; 
      when 1580 => DO <= x"00000000"; 
      when 1581 => DO <= x"00000000"; 
      when 1582 => DO <= x"00000000"; 
      when 1583 => DO <= x"00000000"; 
      when 1584 => DO <= x"00000000"; 
      when 1585 => DO <= x"00000000"; 
      when 1586 => DO <= x"00000000"; 
      when 1587 => DO <= x"00000000"; 
      when 1588 => DO <= x"00000000"; 
      when 1589 => DO <= x"00000000"; 
      when 1590 => DO <= x"00000000"; 
      when 1591 => DO <= x"00000000"; 
      when 1592 => DO <= x"00000000"; 
      when 1593 => DO <= x"00000000"; 
      when 1594 => DO <= x"00000000"; 
      when 1595 => DO <= x"00000000"; 
      when 1596 => DO <= x"00000000"; 
      when 1597 => DO <= x"00000000"; 
      when 1598 => DO <= x"00000000"; 
      when 1599 => DO <= x"00000000"; 
      when 1600 => DO <= x"00000000"; 
      when 1601 => DO <= x"00000000"; 
      when 1602 => DO <= x"00000000"; 
      when 1603 => DO <= x"00000000"; 
      when 1604 => DO <= x"00000000"; 
      when 1605 => DO <= x"00000000"; 
      when 1606 => DO <= x"00000000"; 
      when 1607 => DO <= x"00000000"; 
      when 1608 => DO <= x"00000000"; 
      when 1609 => DO <= x"00000000"; 
      when 1610 => DO <= x"00000000"; 
      when 1611 => DO <= x"00000000"; 
      when 1612 => DO <= x"00000000"; 
      when 1613 => DO <= x"00000000"; 
      when 1614 => DO <= x"00000000"; 
      when 1615 => DO <= x"00000000"; 
      when 1616 => DO <= x"00000000"; 
      when 1617 => DO <= x"00000000"; 
      when 1618 => DO <= x"00000000"; 
      when 1619 => DO <= x"00000000"; 
      when 1620 => DO <= x"00000000"; 
      when 1621 => DO <= x"00000000"; 
      when 1622 => DO <= x"00000000"; 
      when 1623 => DO <= x"00000000"; 
      when 1624 => DO <= x"00000000"; 
      when 1625 => DO <= x"00000000"; 
      when 1626 => DO <= x"00000000"; 
      when 1627 => DO <= x"00000000"; 
      when 1628 => DO <= x"00000000"; 
      when 1629 => DO <= x"00000000"; 
      when 1630 => DO <= x"00000000"; 
      when 1631 => DO <= x"00000000"; 
      when 1632 => DO <= x"00000000"; 
      when 1633 => DO <= x"00000000"; 
      when 1634 => DO <= x"00000000"; 
      when 1635 => DO <= x"00000000"; 
      when 1636 => DO <= x"00000000"; 
      when 1637 => DO <= x"00000000"; 
      when 1638 => DO <= x"00000000"; 
      when 1639 => DO <= x"00000000"; 
      when 1640 => DO <= x"00000000"; 
      when 1641 => DO <= x"00000000"; 
      when 1642 => DO <= x"00000000"; 
      when 1643 => DO <= x"00000000"; 
      when 1644 => DO <= x"00000000"; 
      when 1645 => DO <= x"00000000"; 
      when 1646 => DO <= x"00000000"; 
      when 1647 => DO <= x"00000000"; 
      when 1648 => DO <= x"00000000"; 
      when 1649 => DO <= x"00000000"; 
      when 1650 => DO <= x"00000000"; 
      when 1651 => DO <= x"00000000"; 
      when 1652 => DO <= x"00000000"; 
      when 1653 => DO <= x"00000000"; 
      when 1654 => DO <= x"00000000"; 
      when 1655 => DO <= x"00000000"; 
      when 1656 => DO <= x"00000000"; 
      when 1657 => DO <= x"00000000"; 
      when 1658 => DO <= x"00000000"; 
      when 1659 => DO <= x"00000000"; 
      when 1660 => DO <= x"00000000"; 
      when 1661 => DO <= x"00000000"; 
      when 1662 => DO <= x"00000000"; 
      when 1663 => DO <= x"00000000"; 
      when 1664 => DO <= x"00000000"; 
      when 1665 => DO <= x"00000000"; 
      when 1666 => DO <= x"00000000"; 
      when 1667 => DO <= x"00000000"; 
      when 1668 => DO <= x"00000000"; 
      when 1669 => DO <= x"00000000"; 
      when 1670 => DO <= x"00000000"; 
      when 1671 => DO <= x"00000000"; 
      when 1672 => DO <= x"00000000"; 
      when 1673 => DO <= x"00000000"; 
      when 1674 => DO <= x"00000000"; 
      when 1675 => DO <= x"00000000"; 
      when 1676 => DO <= x"00000000"; 
      when 1677 => DO <= x"00000000"; 
      when 1678 => DO <= x"00000000"; 
      when 1679 => DO <= x"00000000"; 
      when 1680 => DO <= x"00000000"; 
      when 1681 => DO <= x"00000000"; 
      when 1682 => DO <= x"00000000"; 
      when 1683 => DO <= x"00000000"; 
      when 1684 => DO <= x"00000000"; 
      when 1685 => DO <= x"00000000"; 
      when 1686 => DO <= x"00000000"; 
      when 1687 => DO <= x"00000000"; 
      when 1688 => DO <= x"00000000"; 
      when 1689 => DO <= x"00000000"; 
      when 1690 => DO <= x"00000000"; 
      when 1691 => DO <= x"00000000"; 
      when 1692 => DO <= x"00000000"; 
      when 1693 => DO <= x"00000000"; 
      when 1694 => DO <= x"00000000"; 
      when 1695 => DO <= x"00000000"; 
      when 1696 => DO <= x"00000000"; 
      when 1697 => DO <= x"00000000"; 
      when 1698 => DO <= x"00000000"; 
      when 1699 => DO <= x"00000000"; 
      when 1700 => DO <= x"00000000"; 
      when 1701 => DO <= x"00000000"; 
      when 1702 => DO <= x"00000000"; 
      when 1703 => DO <= x"00000000"; 
      when 1704 => DO <= x"00000000"; 
      when 1705 => DO <= x"00000000"; 
      when 1706 => DO <= x"00000000"; 
      when 1707 => DO <= x"00000000"; 
      when 1708 => DO <= x"00000000"; 
      when 1709 => DO <= x"00000000"; 
      when 1710 => DO <= x"00000000"; 
      when 1711 => DO <= x"00000000"; 
      when 1712 => DO <= x"00000000"; 
      when 1713 => DO <= x"00000000"; 
      when 1714 => DO <= x"00000000"; 
      when 1715 => DO <= x"00000000"; 
      when 1716 => DO <= x"00000000"; 
      when 1717 => DO <= x"00000000"; 
      when 1718 => DO <= x"00000000"; 
      when 1719 => DO <= x"00000000"; 
      when 1720 => DO <= x"00000000"; 
      when 1721 => DO <= x"00000000"; 
      when 1722 => DO <= x"00000000"; 
      when 1723 => DO <= x"00000000"; 
      when 1724 => DO <= x"00000000"; 
      when 1725 => DO <= x"00000000"; 
      when 1726 => DO <= x"00000000"; 
      when 1727 => DO <= x"00000000"; 
      when 1728 => DO <= x"00000000"; 
      when 1729 => DO <= x"00000000"; 
      when 1730 => DO <= x"00000000"; 
      when 1731 => DO <= x"00000000"; 
      when 1732 => DO <= x"00000000"; 
      when 1733 => DO <= x"00000000"; 
      when 1734 => DO <= x"00000000"; 
      when 1735 => DO <= x"00000000"; 
      when 1736 => DO <= x"00000000"; 
      when 1737 => DO <= x"00000000"; 
      when 1738 => DO <= x"00000000"; 
      when 1739 => DO <= x"00000000"; 
      when 1740 => DO <= x"00000000"; 
      when 1741 => DO <= x"00000000"; 
      when 1742 => DO <= x"00000000"; 
      when 1743 => DO <= x"00000000"; 
      when 1744 => DO <= x"00000000"; 
      when 1745 => DO <= x"00000000"; 
      when 1746 => DO <= x"00000000"; 
      when 1747 => DO <= x"00000000"; 
      when 1748 => DO <= x"00000000"; 
      when 1749 => DO <= x"00000000"; 
      when 1750 => DO <= x"00000000"; 
      when 1751 => DO <= x"00000000"; 
      when 1752 => DO <= x"00000000"; 
      when 1753 => DO <= x"00000000"; 
      when 1754 => DO <= x"00000000"; 
      when 1755 => DO <= x"00000000"; 
      when 1756 => DO <= x"00000000"; 
      when 1757 => DO <= x"00000000"; 
      when 1758 => DO <= x"00000000"; 
      when 1759 => DO <= x"00000000"; 
      when 1760 => DO <= x"00000000"; 
      when 1761 => DO <= x"00000000"; 
      when 1762 => DO <= x"00000000"; 
      when 1763 => DO <= x"00000000"; 
      when 1764 => DO <= x"00000000"; 
      when 1765 => DO <= x"00000000"; 
      when 1766 => DO <= x"00000000"; 
      when 1767 => DO <= x"00000000"; 
      when 1768 => DO <= x"00000000"; 
      when 1769 => DO <= x"00000000"; 
      when 1770 => DO <= x"00000000"; 
      when 1771 => DO <= x"00000000"; 
      when 1772 => DO <= x"00000000"; 
      when 1773 => DO <= x"00000000"; 
      when 1774 => DO <= x"00000000"; 
      when 1775 => DO <= x"00000000"; 
      when 1776 => DO <= x"00000000"; 
      when 1777 => DO <= x"00000000"; 
      when 1778 => DO <= x"00000000"; 
      when 1779 => DO <= x"00000000"; 
      when 1780 => DO <= x"00000000"; 
      when 1781 => DO <= x"00000000"; 
      when 1782 => DO <= x"00000000"; 
      when 1783 => DO <= x"00000000"; 
      when 1784 => DO <= x"00000000"; 
      when 1785 => DO <= x"00000000"; 
      when 1786 => DO <= x"00000000"; 
      when 1787 => DO <= x"00000000"; 
      when 1788 => DO <= x"00000000"; 
      when 1789 => DO <= x"00000000"; 
      when 1790 => DO <= x"00000000"; 
      when 1791 => DO <= x"00000000"; 
      when 1792 => DO <= x"00000000"; 
      when 1793 => DO <= x"00000000"; 
      when 1794 => DO <= x"00000000"; 
      when 1795 => DO <= x"00000000"; 
      when 1796 => DO <= x"00000000"; 
      when 1797 => DO <= x"00000000"; 
      when 1798 => DO <= x"00000000"; 
      when 1799 => DO <= x"00000000"; 
      when 1800 => DO <= x"00000000"; 
      when 1801 => DO <= x"00000000"; 
      when 1802 => DO <= x"00000000"; 
      when 1803 => DO <= x"00000000"; 
      when 1804 => DO <= x"00000000"; 
      when 1805 => DO <= x"00000000"; 
      when 1806 => DO <= x"00000000"; 
      when 1807 => DO <= x"00000000"; 
      when 1808 => DO <= x"00000000"; 
      when 1809 => DO <= x"00000000"; 
      when 1810 => DO <= x"00000000"; 
      when 1811 => DO <= x"00000000"; 
      when 1812 => DO <= x"00000000"; 
      when 1813 => DO <= x"00000000"; 
      when 1814 => DO <= x"00000000"; 
      when 1815 => DO <= x"00000000"; 
      when 1816 => DO <= x"00000000"; 
      when 1817 => DO <= x"00000000"; 
      when 1818 => DO <= x"00000000"; 
      when 1819 => DO <= x"00000000"; 
      when 1820 => DO <= x"00000000"; 
      when 1821 => DO <= x"00000000"; 
      when 1822 => DO <= x"00000000"; 
      when 1823 => DO <= x"00000000"; 
      when 1824 => DO <= x"00000000"; 
      when 1825 => DO <= x"00000000"; 
      when 1826 => DO <= x"00000000"; 
      when 1827 => DO <= x"00000000"; 
      when 1828 => DO <= x"00000000"; 
      when 1829 => DO <= x"00000000"; 
      when 1830 => DO <= x"00000000"; 
      when 1831 => DO <= x"00000000"; 
      when 1832 => DO <= x"00000000"; 
      when 1833 => DO <= x"00000000"; 
      when 1834 => DO <= x"00000000"; 
      when 1835 => DO <= x"00000000"; 
      when 1836 => DO <= x"00000000"; 
      when 1837 => DO <= x"00000000"; 
      when 1838 => DO <= x"00000000"; 
      when 1839 => DO <= x"00000000"; 
      when 1840 => DO <= x"00000000"; 
      when 1841 => DO <= x"00000000"; 
      when 1842 => DO <= x"00000000"; 
      when 1843 => DO <= x"00000000"; 
      when 1844 => DO <= x"00000000"; 
      when 1845 => DO <= x"00000000"; 
      when 1846 => DO <= x"00000000"; 
      when 1847 => DO <= x"00000000"; 
      when 1848 => DO <= x"00000000"; 
      when 1849 => DO <= x"00000000"; 
      when 1850 => DO <= x"00000000"; 
      when 1851 => DO <= x"00000000"; 
      when 1852 => DO <= x"00000000"; 
      when 1853 => DO <= x"00000000"; 
      when 1854 => DO <= x"00000000"; 
      when 1855 => DO <= x"00000000"; 
      when 1856 => DO <= x"00000000"; 
      when 1857 => DO <= x"00000000"; 
      when 1858 => DO <= x"00000000"; 
      when 1859 => DO <= x"00000000"; 
      when 1860 => DO <= x"00000000"; 
      when 1861 => DO <= x"00000000"; 
      when 1862 => DO <= x"00000000"; 
      when 1863 => DO <= x"00000000"; 
      when 1864 => DO <= x"00000000"; 
      when 1865 => DO <= x"00000000"; 
      when 1866 => DO <= x"00000000"; 
      when 1867 => DO <= x"00000000"; 
      when 1868 => DO <= x"00000000"; 
      when 1869 => DO <= x"00000000"; 
      when 1870 => DO <= x"00000000"; 
      when 1871 => DO <= x"00000000"; 
      when 1872 => DO <= x"00000000"; 
      when 1873 => DO <= x"00000000"; 
      when 1874 => DO <= x"00000000"; 
      when 1875 => DO <= x"00000000"; 
      when 1876 => DO <= x"00000000"; 
      when 1877 => DO <= x"00000000"; 
      when 1878 => DO <= x"00000000"; 
      when 1879 => DO <= x"00000000"; 
      when 1880 => DO <= x"00000000"; 
      when 1881 => DO <= x"00000000"; 
      when 1882 => DO <= x"00000000"; 
      when 1883 => DO <= x"00000000"; 
      when 1884 => DO <= x"00000000"; 
      when 1885 => DO <= x"00000000"; 
      when 1886 => DO <= x"00000000"; 
      when 1887 => DO <= x"00000000"; 
      when 1888 => DO <= x"00000000"; 
      when 1889 => DO <= x"00000000"; 
      when 1890 => DO <= x"00000000"; 
      when 1891 => DO <= x"00000000"; 
      when 1892 => DO <= x"00000000"; 
      when 1893 => DO <= x"00000000"; 
      when 1894 => DO <= x"00000000"; 
      when 1895 => DO <= x"00000000"; 
      when 1896 => DO <= x"00000000"; 
      when 1897 => DO <= x"00000000"; 
      when 1898 => DO <= x"00000000"; 
      when 1899 => DO <= x"00000000"; 
      when 1900 => DO <= x"00000000"; 
      when 1901 => DO <= x"00000000"; 
      when 1902 => DO <= x"00000000"; 
      when 1903 => DO <= x"00000000"; 
      when 1904 => DO <= x"00000000"; 
      when 1905 => DO <= x"00000000"; 
      when 1906 => DO <= x"00000000"; 
      when 1907 => DO <= x"00000000"; 
      when 1908 => DO <= x"00000000"; 
      when 1909 => DO <= x"00000000"; 
      when 1910 => DO <= x"00000000"; 
      when 1911 => DO <= x"00000000"; 
      when 1912 => DO <= x"00000000"; 
      when 1913 => DO <= x"00000000"; 
      when 1914 => DO <= x"00000000"; 
      when 1915 => DO <= x"00000000"; 
      when 1916 => DO <= x"00000000"; 
      when 1917 => DO <= x"00000000"; 
      when 1918 => DO <= x"00000000"; 
      when 1919 => DO <= x"00000000"; 
      when 1920 => DO <= x"00000000"; 
      when 1921 => DO <= x"00000000"; 
      when 1922 => DO <= x"00000000"; 
      when 1923 => DO <= x"00000000"; 
      when 1924 => DO <= x"00000000"; 
      when 1925 => DO <= x"00000000"; 
      when 1926 => DO <= x"00000000"; 
      when 1927 => DO <= x"00000000"; 
      when 1928 => DO <= x"00000000"; 
      when 1929 => DO <= x"00000000"; 
      when 1930 => DO <= x"00000000"; 
      when 1931 => DO <= x"00000000"; 
      when 1932 => DO <= x"00000000"; 
      when 1933 => DO <= x"00000000"; 
      when 1934 => DO <= x"00000000"; 
      when 1935 => DO <= x"00000000"; 
      when 1936 => DO <= x"00000000"; 
      when 1937 => DO <= x"00000000"; 
      when 1938 => DO <= x"00000000"; 
      when 1939 => DO <= x"00000000"; 
      when 1940 => DO <= x"00000000"; 
      when 1941 => DO <= x"00000000"; 
      when 1942 => DO <= x"00000000"; 
      when 1943 => DO <= x"00000000"; 
      when 1944 => DO <= x"00000000"; 
      when 1945 => DO <= x"00000000"; 
      when 1946 => DO <= x"00000000"; 
      when 1947 => DO <= x"00000000"; 
      when 1948 => DO <= x"00000000"; 
      when 1949 => DO <= x"00000000"; 
      when 1950 => DO <= x"00000000"; 
      when 1951 => DO <= x"00000000"; 
      when 1952 => DO <= x"00000000"; 
      when 1953 => DO <= x"00000000"; 
      when 1954 => DO <= x"00000000"; 
      when 1955 => DO <= x"00000000"; 
      when 1956 => DO <= x"00000000"; 
      when 1957 => DO <= x"00000000"; 
      when 1958 => DO <= x"00000000"; 
      when 1959 => DO <= x"00000000"; 
      when 1960 => DO <= x"00000000"; 
      when 1961 => DO <= x"00000000"; 
      when 1962 => DO <= x"00000000"; 
      when 1963 => DO <= x"00000000"; 
      when 1964 => DO <= x"00000000"; 
      when 1965 => DO <= x"00000000"; 
      when 1966 => DO <= x"00000000"; 
      when 1967 => DO <= x"00000000"; 
      when 1968 => DO <= x"00000000"; 
      when 1969 => DO <= x"00000000"; 
      when 1970 => DO <= x"00000000"; 
      when 1971 => DO <= x"00000000"; 
      when 1972 => DO <= x"00000000"; 
      when 1973 => DO <= x"00000000"; 
      when 1974 => DO <= x"00000000"; 
      when 1975 => DO <= x"00000000"; 
      when 1976 => DO <= x"00000000"; 
      when 1977 => DO <= x"00000000"; 
      when 1978 => DO <= x"00000000"; 
      when 1979 => DO <= x"00000000"; 
      when 1980 => DO <= x"00000000"; 
      when 1981 => DO <= x"00000000"; 
      when 1982 => DO <= x"00000000"; 
      when 1983 => DO <= x"00000000"; 
      when 1984 => DO <= x"00000000"; 
      when 1985 => DO <= x"00000000"; 
      when 1986 => DO <= x"00000000"; 
      when 1987 => DO <= x"00000000"; 
      when 1988 => DO <= x"00000000"; 
      when 1989 => DO <= x"00000000"; 
      when 1990 => DO <= x"00000000"; 
      when 1991 => DO <= x"00000000"; 
      when 1992 => DO <= x"00000000"; 
      when 1993 => DO <= x"00000000"; 
      when 1994 => DO <= x"00000000"; 
      when 1995 => DO <= x"00000000"; 
      when 1996 => DO <= x"00000000"; 
      when 1997 => DO <= x"00000000"; 
      when 1998 => DO <= x"00000000"; 
      when 1999 => DO <= x"00000000"; 
      when 2000 => DO <= x"00000000"; 
      when 2001 => DO <= x"00000000"; 
      when 2002 => DO <= x"00000000"; 
      when 2003 => DO <= x"00000000"; 
      when 2004 => DO <= x"00000000"; 
      when 2005 => DO <= x"00000000"; 
      when 2006 => DO <= x"00000000"; 
      when 2007 => DO <= x"00000000"; 
      when 2008 => DO <= x"00000000"; 
      when 2009 => DO <= x"00000000"; 
      when 2010 => DO <= x"00000000"; 
      when 2011 => DO <= x"00000000"; 
      when 2012 => DO <= x"00000000"; 
      when 2013 => DO <= x"00000000"; 
      when 2014 => DO <= x"00000000"; 
      when 2015 => DO <= x"00000000"; 
      when 2016 => DO <= x"00000000"; 
      when 2017 => DO <= x"00000000"; 
      when 2018 => DO <= x"00000000"; 
      when 2019 => DO <= x"00000000"; 
      when 2020 => DO <= x"00000000"; 
      when 2021 => DO <= x"00000000"; 
      when 2022 => DO <= x"00000000"; 
      when 2023 => DO <= x"00000000"; 
      when 2024 => DO <= x"00000000"; 
      when 2025 => DO <= x"00000000"; 
      when 2026 => DO <= x"00000000"; 
      when 2027 => DO <= x"00000000"; 
      when 2028 => DO <= x"00000000"; 
      when 2029 => DO <= x"00000000"; 
      when 2030 => DO <= x"00000000"; 
      when 2031 => DO <= x"00000000"; 
      when 2032 => DO <= x"00000000"; 
      when 2033 => DO <= x"00000000"; 
      when 2034 => DO <= x"00000000"; 
      when 2035 => DO <= x"00000000"; 
      when 2036 => DO <= x"00000000"; 
      when 2037 => DO <= x"00000000"; 
      when 2038 => DO <= x"00000000"; 
      when 2039 => DO <= x"00000000"; 
      when 2040 => DO <= x"00000000"; 
      when 2041 => DO <= x"00000000"; 
      when 2042 => DO <= x"00000000"; 
      when 2043 => DO <= x"00000000"; 
      when 2044 => DO <= x"00000000"; 
      when 2045 => DO <= x"00000000"; 
      when 2046 => DO <= x"00000000"; 
      when 2047 => DO <= x"00000000"; 
when others =>
end case;
end if;
end if;
end process;
end behave;
