library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity internalram is
  port (
    CLK:              in std_logic;
    EN:               in std_logic;
    ADDR:             in std_logic_vector(14 downto 2);
    DO:               out std_logic_vector(31 downto 0)
  );
end entity internalram;

architecture behave of internalram is

begin

process(CLK)
variable iaddr: natural;
begin
  if rising_edge(CLK) then
   if EN='1' then
   iaddr := to_integer(unsigned(ADDR));
     case iaddr is 
      when 0 => DO <= x"81006000"; 
      when 1 => DO <= x"700f8000"; 
      when 2 => DO <= x"70207042"; 
      when 3 => DO <= x"73311012"; 
      when 4 => DO <= x"80017000"; 
      when 5 => DO <= x"70013e31"; 
      when 6 => DO <= x"3c113810"; 
      when 7 => DO <= x"85114010"; 
      when 8 => DO <= x"3e118003"; 
      when 9 => DO <= x"700072c1"; 
      when 10 => DO <= x"41ed3810"; 
      when 11 => DO <= x"c78d4002"; 
      when 12 => DO <= x"38108003"; 
      when 13 => DO <= x"700077b2"; 
      when 14 => DO <= x"60018003"; 
      when 15 => DO <= x"71007722"; 
      when 16 => DO <= x"406d0c21"; 
      when 17 => DO <= x"4fe03810"; 
      when 18 => DO <= x"0c181a18"; 
      when 19 => DO <= x"6001c0e0"; 
      when 20 => DO <= x"42005018"; 
      when 21 => DO <= x"0cd6410d"; 
      when 22 => DO <= x"38100c6d"; 
      when 23 => DO <= x"4ec03810"; 
      when 24 => DO <= x"30d03810"; 
      when 25 => DO <= x"00000000"; 
      when 26 => DO <= x"80007020"; 
      when 27 => DO <= x"70027023"; 
      when 28 => DO <= x"98724004"; 
      when 29 => DO <= x"04376007"; 
      when 30 => DO <= x"cf4041ff"; 
      when 31 => DO <= x"38101012"; 
      when 32 => DO <= x"30d03810"; 
      when 33 => DO <= x"00000000"; 
      when 34 => DO <= x"00008001"; 
      when 35 => DO <= x"7000748d"; 
      when 36 => DO <= x"30d07001"; 
      when 37 => DO <= x"4fe03810"; 
      when 38 => DO <= x"4fe03810"; 
      when 39 => DO <= x"00000000"; 
      when 40 => DO <= x"00000000"; 
      when 41 => DO <= x"00000000"; 
      when 42 => DO <= x"00000000"; 
      when 43 => DO <= x"00000000"; 
      when 44 => DO <= x"00000000"; 
      when 45 => DO <= x"00000000"; 
      when 46 => DO <= x"00000000"; 
      when 47 => DO <= x"00000000"; 
      when 48 => DO <= x"00000000"; 
      when 49 => DO <= x"00000000"; 
      when 50 => DO <= x"00000000"; 
      when 51 => DO <= x"00000000"; 
      when 52 => DO <= x"00000000"; 
      when 53 => DO <= x"00000000"; 
      when 54 => DO <= x"00000000"; 
      when 55 => DO <= x"00000000"; 
      when 56 => DO <= x"00000000"; 
      when 57 => DO <= x"00000000"; 
      when 58 => DO <= x"00000000"; 
      when 59 => DO <= x"00000000"; 
      when 60 => DO <= x"00000000"; 
      when 61 => DO <= x"00000000"; 
      when 62 => DO <= x"00000000"; 
      when 63 => DO <= x"00000000"; 
      when 64 => DO <= x"40203810"; 
      when 65 => DO <= x"3e5ff00f"; 
      when 66 => DO <= x"4010180f"; 
      when 67 => DO <= x"101f902f"; 
      when 68 => DO <= x"40fc903f"; 
      when 69 => DO <= x"40f8904f"; 
      when 70 => DO <= x"40f4905f"; 
      when 71 => DO <= x"40f0906f"; 
      when 72 => DO <= x"40ec907f"; 
      when 73 => DO <= x"40e8908f"; 
      when 74 => DO <= x"40e4909f"; 
      when 75 => DO <= x"40e090af"; 
      when 76 => DO <= x"40dc90bf"; 
      when 77 => DO <= x"40d890cf"; 
      when 78 => DO <= x"40d490df"; 
      when 79 => DO <= x"40d090ef"; 
      when 80 => DO <= x"40cc3c5f"; 
      when 81 => DO <= x"34003810"; 
      when 82 => DO <= x"700130d0"; 
      when 83 => DO <= x"38100000"; 
      when 84 => DO <= x"8911401c"; 
      when 85 => DO <= x"73020521"; 
      when 86 => DO <= x"30d03810"; 
      when 87 => DO <= x"8912401c"; 
      when 88 => DO <= x"73030532"; 
      when 89 => DO <= x"70238000"; 
      when 90 => DO <= x"70209870"; 
      when 91 => DO <= x"40040437"; 
      when 92 => DO <= x"6007cf00"; 
      when 93 => DO <= x"41ff3810"; 
      when 94 => DO <= x"511270f3"; 
      when 95 => DO <= x"80007020"; 
      when 96 => DO <= x"90204000"; 
      when 97 => DO <= x"89124018"; 
      when 98 => DO <= x"04327303"; 
      when 99 => DO <= x"05327023"; 
      when 100 => DO <= x"80007020"; 
      when 101 => DO <= x"98704004"; 
      when 102 => DO <= x"04376007"; 
      when 103 => DO <= x"cf0041ff"; 
      when 104 => DO <= x"38105112"; 
      when 105 => DO <= x"70f38000"; 
      when 106 => DO <= x"70209020"; 
      when 107 => DO <= x"40008912"; 
      when 108 => DO <= x"40140432"; 
      when 109 => DO <= x"73030532"; 
      when 110 => DO <= x"70238000"; 
      when 111 => DO <= x"70209870"; 
      when 112 => DO <= x"40040437"; 
      when 113 => DO <= x"6007cf00"; 
      when 114 => DO <= x"41ff3810"; 
      when 115 => DO <= x"511270f3"; 
      when 116 => DO <= x"80007020"; 
      when 117 => DO <= x"90204000"; 
      when 118 => DO <= x"89124010"; 
      when 119 => DO <= x"04327303"; 
      when 120 => DO <= x"05327023"; 
      when 121 => DO <= x"80007020"; 
      when 122 => DO <= x"98704004"; 
      when 123 => DO <= x"04376007"; 
      when 124 => DO <= x"cf0041ff"; 
      when 125 => DO <= x"38105112"; 
      when 126 => DO <= x"70f38000"; 
      when 127 => DO <= x"70209020"; 
      when 128 => DO <= x"40008912"; 
      when 129 => DO <= x"400c0432"; 
      when 130 => DO <= x"73030532"; 
      when 131 => DO <= x"70238000"; 
      when 132 => DO <= x"70209870"; 
      when 133 => DO <= x"40040437"; 
      when 134 => DO <= x"6007cf00"; 
      when 135 => DO <= x"41ff3810"; 
      when 136 => DO <= x"511270f3"; 
      when 137 => DO <= x"80007020"; 
      when 138 => DO <= x"90204000"; 
      when 139 => DO <= x"89124008"; 
      when 140 => DO <= x"04327303"; 
      when 141 => DO <= x"05327023"; 
      when 142 => DO <= x"80007020"; 
      when 143 => DO <= x"98704004"; 
      when 144 => DO <= x"04376007"; 
      when 145 => DO <= x"cf0041ff"; 
      when 146 => DO <= x"38105112"; 
      when 147 => DO <= x"70f38000"; 
      when 148 => DO <= x"70209020"; 
      when 149 => DO <= x"40008912"; 
      when 150 => DO <= x"40040432"; 
      when 151 => DO <= x"73030532"; 
      when 152 => DO <= x"70238000"; 
      when 153 => DO <= x"70209870"; 
      when 154 => DO <= x"40040437"; 
      when 155 => DO <= x"6007cf00"; 
      when 156 => DO <= x"41ff3810"; 
      when 157 => DO <= x"51128000"; 
      when 158 => DO <= x"70209020"; 
      when 159 => DO <= x"400070f2"; 
      when 160 => DO <= x"04217302"; 
      when 161 => DO <= x"05217022"; 
      when 162 => DO <= x"80007020"; 
      when 163 => DO <= x"98304004"; 
      when 164 => DO <= x"04236003"; 
      when 165 => DO <= x"cf0041ff"; 
      when 166 => DO <= x"38105111"; 
      when 167 => DO <= x"80007020"; 
      when 168 => DO <= x"90104000"; 
      when 169 => DO <= x"30d03810"; 
      when 170 => DO <= x"70028100"; 
      when 171 => DO <= x"60007003"; 
      when 172 => DO <= x"aaaa7055"; 
      when 173 => DO <= x"7aa7fff8"; 
      when 174 => DO <= x"40007209"; 
      when 175 => DO <= x"7201881a"; 
      when 176 => DO <= x"40086001"; 
      when 177 => DO <= x"051a88ab"; 
      when 178 => DO <= x"401005ba"; 
      when 179 => DO <= x"881b4002"; 
      when 180 => DO <= x"067a002b"; 
      when 181 => DO <= x"10ab801a"; 
      when 182 => DO <= x"40ff0ca1"; 
      when 183 => DO <= x"cde041ff"; 
      when 184 => DO <= x"38108489"; 
      when 185 => DO <= x"2001881a"; 
      when 186 => DO <= x"400805a1"; 
      when 187 => DO <= x"881a4010"; 
      when 188 => DO <= x"05a18617"; 
      when 189 => DO <= x"200a8891"; 
      when 190 => DO <= x"40020021"; 
      when 191 => DO <= x"18b17011"; 
      when 192 => DO <= x"07abc200"; 
      when 193 => DO <= x"41003810"; 
      when 194 => DO <= x"809140ff"; 
      when 195 => DO <= x"60090c19"; 
      when 196 => DO <= x"cce041ff"; 
      when 197 => DO <= x"38105ff3"; 
      when 198 => DO <= x"d8024000"; 
      when 199 => DO <= x"70016003"; 
      when 200 => DO <= x"c96041ff"; 
      when 201 => DO <= x"381030d0"; 
      when 202 => DO <= x"38100000"; 
      when 203 => DO <= x"58546875"; 
      when 204 => DO <= x"6e646572"; 
      when 205 => DO <= x"436f7265"; 
      when 206 => DO <= x"20426f6f"; 
      when 207 => DO <= x"74204c6f"; 
      when 208 => DO <= x"61646572"; 
      when 209 => DO <= x"2076302e"; 
      when 210 => DO <= x"31202843"; 
      when 211 => DO <= x"29203230"; 
      when 212 => DO <= x"31342041"; 
      when 213 => DO <= x"6c766172"; 
      when 214 => DO <= x"6f204c6f"; 
      when 215 => DO <= x"7065730d"; 
      when 216 => DO <= x"0a546573"; 
      when 217 => DO <= x"74696e67"; 
      when 218 => DO <= x"206d656d"; 
      when 219 => DO <= x"6f72793a"; 
      when 220 => DO <= x"20004661"; 
      when 221 => DO <= x"696c6564"; 
      when 222 => DO <= x"0d0a0050"; 
      when 223 => DO <= x"61737365"; 
      when 224 => DO <= x"640d0a00"; 
      when 225 => DO <= x"00000000"; 
      when 226 => DO <= x"00000000"; 
      when 227 => DO <= x"00000000"; 
      when 228 => DO <= x"00000000"; 
      when 229 => DO <= x"00000000"; 
      when 230 => DO <= x"00000000"; 
      when 231 => DO <= x"00000000"; 
      when 232 => DO <= x"00000000"; 
      when 233 => DO <= x"00000000"; 
      when 234 => DO <= x"00000000"; 
      when 235 => DO <= x"00000000"; 
      when 236 => DO <= x"00000000"; 
      when 237 => DO <= x"00000000"; 
      when 238 => DO <= x"00000000"; 
      when 239 => DO <= x"00000000"; 
      when 240 => DO <= x"00000000"; 
      when 241 => DO <= x"00000000"; 
      when 242 => DO <= x"00000000"; 
      when 243 => DO <= x"00000000"; 
      when 244 => DO <= x"00000000"; 
      when 245 => DO <= x"00000000"; 
      when 246 => DO <= x"00000000"; 
      when 247 => DO <= x"00000000"; 
      when 248 => DO <= x"00000000"; 
      when 249 => DO <= x"00000000"; 
      when 250 => DO <= x"00000000"; 
      when 251 => DO <= x"00000000"; 
      when 252 => DO <= x"00000000"; 
      when 253 => DO <= x"00000000"; 
      when 254 => DO <= x"00000000"; 
      when 255 => DO <= x"00000000"; 
      when 256 => DO <= x"00000000"; 
      when 257 => DO <= x"00000000"; 
      when 258 => DO <= x"00000000"; 
      when 259 => DO <= x"00000000"; 
      when 260 => DO <= x"00000000"; 
      when 261 => DO <= x"00000000"; 
      when 262 => DO <= x"00000000"; 
      when 263 => DO <= x"00000000"; 
      when 264 => DO <= x"00000000"; 
      when 265 => DO <= x"00000000"; 
      when 266 => DO <= x"00000000"; 
      when 267 => DO <= x"00000000"; 
      when 268 => DO <= x"00000000"; 
      when 269 => DO <= x"00000000"; 
      when 270 => DO <= x"00000000"; 
      when 271 => DO <= x"00000000"; 
      when 272 => DO <= x"00000000"; 
      when 273 => DO <= x"00000000"; 
      when 274 => DO <= x"00000000"; 
      when 275 => DO <= x"00000000"; 
      when 276 => DO <= x"00000000"; 
      when 277 => DO <= x"00000000"; 
      when 278 => DO <= x"00000000"; 
      when 279 => DO <= x"00000000"; 
      when 280 => DO <= x"00000000"; 
      when 281 => DO <= x"00000000"; 
      when 282 => DO <= x"00000000"; 
      when 283 => DO <= x"00000000"; 
      when 284 => DO <= x"00000000"; 
      when 285 => DO <= x"00000000"; 
      when 286 => DO <= x"00000000"; 
      when 287 => DO <= x"00000000"; 
      when 288 => DO <= x"00000000"; 
      when 289 => DO <= x"00000000"; 
      when 290 => DO <= x"00000000"; 
      when 291 => DO <= x"00000000"; 
      when 292 => DO <= x"00000000"; 
      when 293 => DO <= x"00000000"; 
      when 294 => DO <= x"00000000"; 
      when 295 => DO <= x"00000000"; 
      when 296 => DO <= x"00000000"; 
      when 297 => DO <= x"00000000"; 
      when 298 => DO <= x"00000000"; 
      when 299 => DO <= x"00000000"; 
      when 300 => DO <= x"00000000"; 
      when 301 => DO <= x"00000000"; 
      when 302 => DO <= x"00000000"; 
      when 303 => DO <= x"00000000"; 
      when 304 => DO <= x"00000000"; 
      when 305 => DO <= x"00000000"; 
      when 306 => DO <= x"00000000"; 
      when 307 => DO <= x"00000000"; 
      when 308 => DO <= x"00000000"; 
      when 309 => DO <= x"00000000"; 
      when 310 => DO <= x"00000000"; 
      when 311 => DO <= x"00000000"; 
      when 312 => DO <= x"00000000"; 
      when 313 => DO <= x"00000000"; 
      when 314 => DO <= x"00000000"; 
      when 315 => DO <= x"00000000"; 
      when 316 => DO <= x"00000000"; 
      when 317 => DO <= x"00000000"; 
      when 318 => DO <= x"00000000"; 
      when 319 => DO <= x"00000000"; 
      when 320 => DO <= x"00000000"; 
      when 321 => DO <= x"00000000"; 
      when 322 => DO <= x"00000000"; 
      when 323 => DO <= x"00000000"; 
      when 324 => DO <= x"00000000"; 
      when 325 => DO <= x"00000000"; 
      when 326 => DO <= x"00000000"; 
      when 327 => DO <= x"00000000"; 
      when 328 => DO <= x"00000000"; 
      when 329 => DO <= x"00000000"; 
      when 330 => DO <= x"00000000"; 
      when 331 => DO <= x"00000000"; 
      when 332 => DO <= x"00000000"; 
      when 333 => DO <= x"00000000"; 
      when 334 => DO <= x"00000000"; 
      when 335 => DO <= x"00000000"; 
      when 336 => DO <= x"00000000"; 
      when 337 => DO <= x"00000000"; 
      when 338 => DO <= x"00000000"; 
      when 339 => DO <= x"00000000"; 
      when 340 => DO <= x"00000000"; 
      when 341 => DO <= x"00000000"; 
      when 342 => DO <= x"00000000"; 
      when 343 => DO <= x"00000000"; 
      when 344 => DO <= x"00000000"; 
      when 345 => DO <= x"00000000"; 
      when 346 => DO <= x"00000000"; 
      when 347 => DO <= x"00000000"; 
      when 348 => DO <= x"00000000"; 
      when 349 => DO <= x"00000000"; 
      when 350 => DO <= x"00000000"; 
      when 351 => DO <= x"00000000"; 
      when 352 => DO <= x"00000000"; 
      when 353 => DO <= x"00000000"; 
      when 354 => DO <= x"00000000"; 
      when 355 => DO <= x"00000000"; 
      when 356 => DO <= x"00000000"; 
      when 357 => DO <= x"00000000"; 
      when 358 => DO <= x"00000000"; 
      when 359 => DO <= x"00000000"; 
      when 360 => DO <= x"00000000"; 
      when 361 => DO <= x"00000000"; 
      when 362 => DO <= x"00000000"; 
      when 363 => DO <= x"00000000"; 
      when 364 => DO <= x"00000000"; 
      when 365 => DO <= x"00000000"; 
      when 366 => DO <= x"00000000"; 
      when 367 => DO <= x"00000000"; 
      when 368 => DO <= x"00000000"; 
      when 369 => DO <= x"00000000"; 
      when 370 => DO <= x"00000000"; 
      when 371 => DO <= x"00000000"; 
      when 372 => DO <= x"00000000"; 
      when 373 => DO <= x"00000000"; 
      when 374 => DO <= x"00000000"; 
      when 375 => DO <= x"00000000"; 
      when 376 => DO <= x"00000000"; 
      when 377 => DO <= x"00000000"; 
      when 378 => DO <= x"00000000"; 
      when 379 => DO <= x"00000000"; 
      when 380 => DO <= x"00000000"; 
      when 381 => DO <= x"00000000"; 
      when 382 => DO <= x"00000000"; 
      when 383 => DO <= x"00000000"; 
      when 384 => DO <= x"00000000"; 
      when 385 => DO <= x"00000000"; 
      when 386 => DO <= x"00000000"; 
      when 387 => DO <= x"00000000"; 
      when 388 => DO <= x"00000000"; 
      when 389 => DO <= x"00000000"; 
      when 390 => DO <= x"00000000"; 
      when 391 => DO <= x"00000000"; 
      when 392 => DO <= x"00000000"; 
      when 393 => DO <= x"00000000"; 
      when 394 => DO <= x"00000000"; 
      when 395 => DO <= x"00000000"; 
      when 396 => DO <= x"00000000"; 
      when 397 => DO <= x"00000000"; 
      when 398 => DO <= x"00000000"; 
      when 399 => DO <= x"00000000"; 
      when 400 => DO <= x"00000000"; 
      when 401 => DO <= x"00000000"; 
      when 402 => DO <= x"00000000"; 
      when 403 => DO <= x"00000000"; 
      when 404 => DO <= x"00000000"; 
      when 405 => DO <= x"00000000"; 
      when 406 => DO <= x"00000000"; 
      when 407 => DO <= x"00000000"; 
      when 408 => DO <= x"00000000"; 
      when 409 => DO <= x"00000000"; 
      when 410 => DO <= x"00000000"; 
      when 411 => DO <= x"00000000"; 
      when 412 => DO <= x"00000000"; 
      when 413 => DO <= x"00000000"; 
      when 414 => DO <= x"00000000"; 
      when 415 => DO <= x"00000000"; 
      when 416 => DO <= x"00000000"; 
      when 417 => DO <= x"00000000"; 
      when 418 => DO <= x"00000000"; 
      when 419 => DO <= x"00000000"; 
      when 420 => DO <= x"00000000"; 
      when 421 => DO <= x"00000000"; 
      when 422 => DO <= x"00000000"; 
      when 423 => DO <= x"00000000"; 
      when 424 => DO <= x"00000000"; 
      when 425 => DO <= x"00000000"; 
      when 426 => DO <= x"00000000"; 
      when 427 => DO <= x"00000000"; 
      when 428 => DO <= x"00000000"; 
      when 429 => DO <= x"00000000"; 
      when 430 => DO <= x"00000000"; 
      when 431 => DO <= x"00000000"; 
      when 432 => DO <= x"00000000"; 
      when 433 => DO <= x"00000000"; 
      when 434 => DO <= x"00000000"; 
      when 435 => DO <= x"00000000"; 
      when 436 => DO <= x"00000000"; 
      when 437 => DO <= x"00000000"; 
      when 438 => DO <= x"00000000"; 
      when 439 => DO <= x"00000000"; 
      when 440 => DO <= x"00000000"; 
      when 441 => DO <= x"00000000"; 
      when 442 => DO <= x"00000000"; 
      when 443 => DO <= x"00000000"; 
      when 444 => DO <= x"00000000"; 
      when 445 => DO <= x"00000000"; 
      when 446 => DO <= x"00000000"; 
      when 447 => DO <= x"00000000"; 
      when 448 => DO <= x"00000000"; 
      when 449 => DO <= x"00000000"; 
      when 450 => DO <= x"00000000"; 
      when 451 => DO <= x"00000000"; 
      when 452 => DO <= x"00000000"; 
      when 453 => DO <= x"00000000"; 
      when 454 => DO <= x"00000000"; 
      when 455 => DO <= x"00000000"; 
      when 456 => DO <= x"00000000"; 
      when 457 => DO <= x"00000000"; 
      when 458 => DO <= x"00000000"; 
      when 459 => DO <= x"00000000"; 
      when 460 => DO <= x"00000000"; 
      when 461 => DO <= x"00000000"; 
      when 462 => DO <= x"00000000"; 
      when 463 => DO <= x"00000000"; 
      when 464 => DO <= x"00000000"; 
      when 465 => DO <= x"00000000"; 
      when 466 => DO <= x"00000000"; 
      when 467 => DO <= x"00000000"; 
      when 468 => DO <= x"00000000"; 
      when 469 => DO <= x"00000000"; 
      when 470 => DO <= x"00000000"; 
      when 471 => DO <= x"00000000"; 
      when 472 => DO <= x"00000000"; 
      when 473 => DO <= x"00000000"; 
      when 474 => DO <= x"00000000"; 
      when 475 => DO <= x"00000000"; 
      when 476 => DO <= x"00000000"; 
      when 477 => DO <= x"00000000"; 
      when 478 => DO <= x"00000000"; 
      when 479 => DO <= x"00000000"; 
      when 480 => DO <= x"00000000"; 
      when 481 => DO <= x"00000000"; 
      when 482 => DO <= x"00000000"; 
      when 483 => DO <= x"00000000"; 
      when 484 => DO <= x"00000000"; 
      when 485 => DO <= x"00000000"; 
      when 486 => DO <= x"00000000"; 
      when 487 => DO <= x"00000000"; 
      when 488 => DO <= x"00000000"; 
      when 489 => DO <= x"00000000"; 
      when 490 => DO <= x"00000000"; 
      when 491 => DO <= x"00000000"; 
      when 492 => DO <= x"00000000"; 
      when 493 => DO <= x"00000000"; 
      when 494 => DO <= x"00000000"; 
      when 495 => DO <= x"00000000"; 
      when 496 => DO <= x"00000000"; 
      when 497 => DO <= x"00000000"; 
      when 498 => DO <= x"00000000"; 
      when 499 => DO <= x"00000000"; 
      when 500 => DO <= x"00000000"; 
      when 501 => DO <= x"00000000"; 
      when 502 => DO <= x"00000000"; 
      when 503 => DO <= x"00000000"; 
      when 504 => DO <= x"00000000"; 
      when 505 => DO <= x"00000000"; 
      when 506 => DO <= x"00000000"; 
      when 507 => DO <= x"00000000"; 
      when 508 => DO <= x"00000000"; 
      when 509 => DO <= x"00000000"; 
      when 510 => DO <= x"00000000"; 
      when 511 => DO <= x"00000000"; 
      when 512 => DO <= x"00000000"; 
      when 513 => DO <= x"00000000"; 
      when 514 => DO <= x"00000000"; 
      when 515 => DO <= x"00000000"; 
      when 516 => DO <= x"00000000"; 
      when 517 => DO <= x"00000000"; 
      when 518 => DO <= x"00000000"; 
      when 519 => DO <= x"00000000"; 
      when 520 => DO <= x"00000000"; 
      when 521 => DO <= x"00000000"; 
      when 522 => DO <= x"00000000"; 
      when 523 => DO <= x"00000000"; 
      when 524 => DO <= x"00000000"; 
      when 525 => DO <= x"00000000"; 
      when 526 => DO <= x"00000000"; 
      when 527 => DO <= x"00000000"; 
      when 528 => DO <= x"00000000"; 
      when 529 => DO <= x"00000000"; 
      when 530 => DO <= x"00000000"; 
      when 531 => DO <= x"00000000"; 
      when 532 => DO <= x"00000000"; 
      when 533 => DO <= x"00000000"; 
      when 534 => DO <= x"00000000"; 
      when 535 => DO <= x"00000000"; 
      when 536 => DO <= x"00000000"; 
      when 537 => DO <= x"00000000"; 
      when 538 => DO <= x"00000000"; 
      when 539 => DO <= x"00000000"; 
      when 540 => DO <= x"00000000"; 
      when 541 => DO <= x"00000000"; 
      when 542 => DO <= x"00000000"; 
      when 543 => DO <= x"00000000"; 
      when 544 => DO <= x"00000000"; 
      when 545 => DO <= x"00000000"; 
      when 546 => DO <= x"00000000"; 
      when 547 => DO <= x"00000000"; 
      when 548 => DO <= x"00000000"; 
      when 549 => DO <= x"00000000"; 
      when 550 => DO <= x"00000000"; 
      when 551 => DO <= x"00000000"; 
      when 552 => DO <= x"00000000"; 
      when 553 => DO <= x"00000000"; 
      when 554 => DO <= x"00000000"; 
      when 555 => DO <= x"00000000"; 
      when 556 => DO <= x"00000000"; 
      when 557 => DO <= x"00000000"; 
      when 558 => DO <= x"00000000"; 
      when 559 => DO <= x"00000000"; 
      when 560 => DO <= x"00000000"; 
      when 561 => DO <= x"00000000"; 
      when 562 => DO <= x"00000000"; 
      when 563 => DO <= x"00000000"; 
      when 564 => DO <= x"00000000"; 
      when 565 => DO <= x"00000000"; 
      when 566 => DO <= x"00000000"; 
      when 567 => DO <= x"00000000"; 
      when 568 => DO <= x"00000000"; 
      when 569 => DO <= x"00000000"; 
      when 570 => DO <= x"00000000"; 
      when 571 => DO <= x"00000000"; 
      when 572 => DO <= x"00000000"; 
      when 573 => DO <= x"00000000"; 
      when 574 => DO <= x"00000000"; 
      when 575 => DO <= x"00000000"; 
      when 576 => DO <= x"00000000"; 
      when 577 => DO <= x"00000000"; 
      when 578 => DO <= x"00000000"; 
      when 579 => DO <= x"00000000"; 
      when 580 => DO <= x"00000000"; 
      when 581 => DO <= x"00000000"; 
      when 582 => DO <= x"00000000"; 
      when 583 => DO <= x"00000000"; 
      when 584 => DO <= x"00000000"; 
      when 585 => DO <= x"00000000"; 
      when 586 => DO <= x"00000000"; 
      when 587 => DO <= x"00000000"; 
      when 588 => DO <= x"00000000"; 
      when 589 => DO <= x"00000000"; 
      when 590 => DO <= x"00000000"; 
      when 591 => DO <= x"00000000"; 
      when 592 => DO <= x"00000000"; 
      when 593 => DO <= x"00000000"; 
      when 594 => DO <= x"00000000"; 
      when 595 => DO <= x"00000000"; 
      when 596 => DO <= x"00000000"; 
      when 597 => DO <= x"00000000"; 
      when 598 => DO <= x"00000000"; 
      when 599 => DO <= x"00000000"; 
      when 600 => DO <= x"00000000"; 
      when 601 => DO <= x"00000000"; 
      when 602 => DO <= x"00000000"; 
      when 603 => DO <= x"00000000"; 
      when 604 => DO <= x"00000000"; 
      when 605 => DO <= x"00000000"; 
      when 606 => DO <= x"00000000"; 
      when 607 => DO <= x"00000000"; 
      when 608 => DO <= x"00000000"; 
      when 609 => DO <= x"00000000"; 
      when 610 => DO <= x"00000000"; 
      when 611 => DO <= x"00000000"; 
      when 612 => DO <= x"00000000"; 
      when 613 => DO <= x"00000000"; 
      when 614 => DO <= x"00000000"; 
      when 615 => DO <= x"00000000"; 
      when 616 => DO <= x"00000000"; 
      when 617 => DO <= x"00000000"; 
      when 618 => DO <= x"00000000"; 
      when 619 => DO <= x"00000000"; 
      when 620 => DO <= x"00000000"; 
      when 621 => DO <= x"00000000"; 
      when 622 => DO <= x"00000000"; 
      when 623 => DO <= x"00000000"; 
      when 624 => DO <= x"00000000"; 
      when 625 => DO <= x"00000000"; 
      when 626 => DO <= x"00000000"; 
      when 627 => DO <= x"00000000"; 
      when 628 => DO <= x"00000000"; 
      when 629 => DO <= x"00000000"; 
      when 630 => DO <= x"00000000"; 
      when 631 => DO <= x"00000000"; 
      when 632 => DO <= x"00000000"; 
      when 633 => DO <= x"00000000"; 
      when 634 => DO <= x"00000000"; 
      when 635 => DO <= x"00000000"; 
      when 636 => DO <= x"00000000"; 
      when 637 => DO <= x"00000000"; 
      when 638 => DO <= x"00000000"; 
      when 639 => DO <= x"00000000"; 
      when 640 => DO <= x"00000000"; 
      when 641 => DO <= x"00000000"; 
      when 642 => DO <= x"00000000"; 
      when 643 => DO <= x"00000000"; 
      when 644 => DO <= x"00000000"; 
      when 645 => DO <= x"00000000"; 
      when 646 => DO <= x"00000000"; 
      when 647 => DO <= x"00000000"; 
      when 648 => DO <= x"00000000"; 
      when 649 => DO <= x"00000000"; 
      when 650 => DO <= x"00000000"; 
      when 651 => DO <= x"00000000"; 
      when 652 => DO <= x"00000000"; 
      when 653 => DO <= x"00000000"; 
      when 654 => DO <= x"00000000"; 
      when 655 => DO <= x"00000000"; 
      when 656 => DO <= x"00000000"; 
      when 657 => DO <= x"00000000"; 
      when 658 => DO <= x"00000000"; 
      when 659 => DO <= x"00000000"; 
      when 660 => DO <= x"00000000"; 
      when 661 => DO <= x"00000000"; 
      when 662 => DO <= x"00000000"; 
      when 663 => DO <= x"00000000"; 
      when 664 => DO <= x"00000000"; 
      when 665 => DO <= x"00000000"; 
      when 666 => DO <= x"00000000"; 
      when 667 => DO <= x"00000000"; 
      when 668 => DO <= x"00000000"; 
      when 669 => DO <= x"00000000"; 
      when 670 => DO <= x"00000000"; 
      when 671 => DO <= x"00000000"; 
      when 672 => DO <= x"00000000"; 
      when 673 => DO <= x"00000000"; 
      when 674 => DO <= x"00000000"; 
      when 675 => DO <= x"00000000"; 
      when 676 => DO <= x"00000000"; 
      when 677 => DO <= x"00000000"; 
      when 678 => DO <= x"00000000"; 
      when 679 => DO <= x"00000000"; 
      when 680 => DO <= x"00000000"; 
      when 681 => DO <= x"00000000"; 
      when 682 => DO <= x"00000000"; 
      when 683 => DO <= x"00000000"; 
      when 684 => DO <= x"00000000"; 
      when 685 => DO <= x"00000000"; 
      when 686 => DO <= x"00000000"; 
      when 687 => DO <= x"00000000"; 
      when 688 => DO <= x"00000000"; 
      when 689 => DO <= x"00000000"; 
      when 690 => DO <= x"00000000"; 
      when 691 => DO <= x"00000000"; 
      when 692 => DO <= x"00000000"; 
      when 693 => DO <= x"00000000"; 
      when 694 => DO <= x"00000000"; 
      when 695 => DO <= x"00000000"; 
      when 696 => DO <= x"00000000"; 
      when 697 => DO <= x"00000000"; 
      when 698 => DO <= x"00000000"; 
      when 699 => DO <= x"00000000"; 
      when 700 => DO <= x"00000000"; 
      when 701 => DO <= x"00000000"; 
      when 702 => DO <= x"00000000"; 
      when 703 => DO <= x"00000000"; 
      when 704 => DO <= x"00000000"; 
      when 705 => DO <= x"00000000"; 
      when 706 => DO <= x"00000000"; 
      when 707 => DO <= x"00000000"; 
      when 708 => DO <= x"00000000"; 
      when 709 => DO <= x"00000000"; 
      when 710 => DO <= x"00000000"; 
      when 711 => DO <= x"00000000"; 
      when 712 => DO <= x"00000000"; 
      when 713 => DO <= x"00000000"; 
      when 714 => DO <= x"00000000"; 
      when 715 => DO <= x"00000000"; 
      when 716 => DO <= x"00000000"; 
      when 717 => DO <= x"00000000"; 
      when 718 => DO <= x"00000000"; 
      when 719 => DO <= x"00000000"; 
      when 720 => DO <= x"00000000"; 
      when 721 => DO <= x"00000000"; 
      when 722 => DO <= x"00000000"; 
      when 723 => DO <= x"00000000"; 
      when 724 => DO <= x"00000000"; 
      when 725 => DO <= x"00000000"; 
      when 726 => DO <= x"00000000"; 
      when 727 => DO <= x"00000000"; 
      when 728 => DO <= x"00000000"; 
      when 729 => DO <= x"00000000"; 
      when 730 => DO <= x"00000000"; 
      when 731 => DO <= x"00000000"; 
      when 732 => DO <= x"00000000"; 
      when 733 => DO <= x"00000000"; 
      when 734 => DO <= x"00000000"; 
      when 735 => DO <= x"00000000"; 
      when 736 => DO <= x"00000000"; 
      when 737 => DO <= x"00000000"; 
      when 738 => DO <= x"00000000"; 
      when 739 => DO <= x"00000000"; 
      when 740 => DO <= x"00000000"; 
      when 741 => DO <= x"00000000"; 
      when 742 => DO <= x"00000000"; 
      when 743 => DO <= x"00000000"; 
      when 744 => DO <= x"00000000"; 
      when 745 => DO <= x"00000000"; 
      when 746 => DO <= x"00000000"; 
      when 747 => DO <= x"00000000"; 
      when 748 => DO <= x"00000000"; 
      when 749 => DO <= x"00000000"; 
      when 750 => DO <= x"00000000"; 
      when 751 => DO <= x"00000000"; 
      when 752 => DO <= x"00000000"; 
      when 753 => DO <= x"00000000"; 
      when 754 => DO <= x"00000000"; 
      when 755 => DO <= x"00000000"; 
      when 756 => DO <= x"00000000"; 
      when 757 => DO <= x"00000000"; 
      when 758 => DO <= x"00000000"; 
      when 759 => DO <= x"00000000"; 
      when 760 => DO <= x"00000000"; 
      when 761 => DO <= x"00000000"; 
      when 762 => DO <= x"00000000"; 
      when 763 => DO <= x"00000000"; 
      when 764 => DO <= x"00000000"; 
      when 765 => DO <= x"00000000"; 
      when 766 => DO <= x"00000000"; 
      when 767 => DO <= x"00000000"; 
      when 768 => DO <= x"00000000"; 
      when 769 => DO <= x"00000000"; 
      when 770 => DO <= x"00000000"; 
      when 771 => DO <= x"00000000"; 
      when 772 => DO <= x"00000000"; 
      when 773 => DO <= x"00000000"; 
      when 774 => DO <= x"00000000"; 
      when 775 => DO <= x"00000000"; 
      when 776 => DO <= x"00000000"; 
      when 777 => DO <= x"00000000"; 
      when 778 => DO <= x"00000000"; 
      when 779 => DO <= x"00000000"; 
      when 780 => DO <= x"00000000"; 
      when 781 => DO <= x"00000000"; 
      when 782 => DO <= x"00000000"; 
      when 783 => DO <= x"00000000"; 
      when 784 => DO <= x"00000000"; 
      when 785 => DO <= x"00000000"; 
      when 786 => DO <= x"00000000"; 
      when 787 => DO <= x"00000000"; 
      when 788 => DO <= x"00000000"; 
      when 789 => DO <= x"00000000"; 
      when 790 => DO <= x"00000000"; 
      when 791 => DO <= x"00000000"; 
      when 792 => DO <= x"00000000"; 
      when 793 => DO <= x"00000000"; 
      when 794 => DO <= x"00000000"; 
      when 795 => DO <= x"00000000"; 
      when 796 => DO <= x"00000000"; 
      when 797 => DO <= x"00000000"; 
      when 798 => DO <= x"00000000"; 
      when 799 => DO <= x"00000000"; 
      when 800 => DO <= x"00000000"; 
      when 801 => DO <= x"00000000"; 
      when 802 => DO <= x"00000000"; 
      when 803 => DO <= x"00000000"; 
      when 804 => DO <= x"00000000"; 
      when 805 => DO <= x"00000000"; 
      when 806 => DO <= x"00000000"; 
      when 807 => DO <= x"00000000"; 
      when 808 => DO <= x"00000000"; 
      when 809 => DO <= x"00000000"; 
      when 810 => DO <= x"00000000"; 
      when 811 => DO <= x"00000000"; 
      when 812 => DO <= x"00000000"; 
      when 813 => DO <= x"00000000"; 
      when 814 => DO <= x"00000000"; 
      when 815 => DO <= x"00000000"; 
      when 816 => DO <= x"00000000"; 
      when 817 => DO <= x"00000000"; 
      when 818 => DO <= x"00000000"; 
      when 819 => DO <= x"00000000"; 
      when 820 => DO <= x"00000000"; 
      when 821 => DO <= x"00000000"; 
      when 822 => DO <= x"00000000"; 
      when 823 => DO <= x"00000000"; 
      when 824 => DO <= x"00000000"; 
      when 825 => DO <= x"00000000"; 
      when 826 => DO <= x"00000000"; 
      when 827 => DO <= x"00000000"; 
      when 828 => DO <= x"00000000"; 
      when 829 => DO <= x"00000000"; 
      when 830 => DO <= x"00000000"; 
      when 831 => DO <= x"00000000"; 
      when 832 => DO <= x"00000000"; 
      when 833 => DO <= x"00000000"; 
      when 834 => DO <= x"00000000"; 
      when 835 => DO <= x"00000000"; 
      when 836 => DO <= x"00000000"; 
      when 837 => DO <= x"00000000"; 
      when 838 => DO <= x"00000000"; 
      when 839 => DO <= x"00000000"; 
      when 840 => DO <= x"00000000"; 
      when 841 => DO <= x"00000000"; 
      when 842 => DO <= x"00000000"; 
      when 843 => DO <= x"00000000"; 
      when 844 => DO <= x"00000000"; 
      when 845 => DO <= x"00000000"; 
      when 846 => DO <= x"00000000"; 
      when 847 => DO <= x"00000000"; 
      when 848 => DO <= x"00000000"; 
      when 849 => DO <= x"00000000"; 
      when 850 => DO <= x"00000000"; 
      when 851 => DO <= x"00000000"; 
      when 852 => DO <= x"00000000"; 
      when 853 => DO <= x"00000000"; 
      when 854 => DO <= x"00000000"; 
      when 855 => DO <= x"00000000"; 
      when 856 => DO <= x"00000000"; 
      when 857 => DO <= x"00000000"; 
      when 858 => DO <= x"00000000"; 
      when 859 => DO <= x"00000000"; 
      when 860 => DO <= x"00000000"; 
      when 861 => DO <= x"00000000"; 
      when 862 => DO <= x"00000000"; 
      when 863 => DO <= x"00000000"; 
      when 864 => DO <= x"00000000"; 
      when 865 => DO <= x"00000000"; 
      when 866 => DO <= x"00000000"; 
      when 867 => DO <= x"00000000"; 
      when 868 => DO <= x"00000000"; 
      when 869 => DO <= x"00000000"; 
      when 870 => DO <= x"00000000"; 
      when 871 => DO <= x"00000000"; 
      when 872 => DO <= x"00000000"; 
      when 873 => DO <= x"00000000"; 
      when 874 => DO <= x"00000000"; 
      when 875 => DO <= x"00000000"; 
      when 876 => DO <= x"00000000"; 
      when 877 => DO <= x"00000000"; 
      when 878 => DO <= x"00000000"; 
      when 879 => DO <= x"00000000"; 
      when 880 => DO <= x"00000000"; 
      when 881 => DO <= x"00000000"; 
      when 882 => DO <= x"00000000"; 
      when 883 => DO <= x"00000000"; 
      when 884 => DO <= x"00000000"; 
      when 885 => DO <= x"00000000"; 
      when 886 => DO <= x"00000000"; 
      when 887 => DO <= x"00000000"; 
      when 888 => DO <= x"00000000"; 
      when 889 => DO <= x"00000000"; 
      when 890 => DO <= x"00000000"; 
      when 891 => DO <= x"00000000"; 
      when 892 => DO <= x"00000000"; 
      when 893 => DO <= x"00000000"; 
      when 894 => DO <= x"00000000"; 
      when 895 => DO <= x"00000000"; 
      when 896 => DO <= x"00000000"; 
      when 897 => DO <= x"00000000"; 
      when 898 => DO <= x"00000000"; 
      when 899 => DO <= x"00000000"; 
      when 900 => DO <= x"00000000"; 
      when 901 => DO <= x"00000000"; 
      when 902 => DO <= x"00000000"; 
      when 903 => DO <= x"00000000"; 
      when 904 => DO <= x"00000000"; 
      when 905 => DO <= x"00000000"; 
      when 906 => DO <= x"00000000"; 
      when 907 => DO <= x"00000000"; 
      when 908 => DO <= x"00000000"; 
      when 909 => DO <= x"00000000"; 
      when 910 => DO <= x"00000000"; 
      when 911 => DO <= x"00000000"; 
      when 912 => DO <= x"00000000"; 
      when 913 => DO <= x"00000000"; 
      when 914 => DO <= x"00000000"; 
      when 915 => DO <= x"00000000"; 
      when 916 => DO <= x"00000000"; 
      when 917 => DO <= x"00000000"; 
      when 918 => DO <= x"00000000"; 
      when 919 => DO <= x"00000000"; 
      when 920 => DO <= x"00000000"; 
      when 921 => DO <= x"00000000"; 
      when 922 => DO <= x"00000000"; 
      when 923 => DO <= x"00000000"; 
      when 924 => DO <= x"00000000"; 
      when 925 => DO <= x"00000000"; 
      when 926 => DO <= x"00000000"; 
      when 927 => DO <= x"00000000"; 
      when 928 => DO <= x"00000000"; 
      when 929 => DO <= x"00000000"; 
      when 930 => DO <= x"00000000"; 
      when 931 => DO <= x"00000000"; 
      when 932 => DO <= x"00000000"; 
      when 933 => DO <= x"00000000"; 
      when 934 => DO <= x"00000000"; 
      when 935 => DO <= x"00000000"; 
      when 936 => DO <= x"00000000"; 
      when 937 => DO <= x"00000000"; 
      when 938 => DO <= x"00000000"; 
      when 939 => DO <= x"00000000"; 
      when 940 => DO <= x"00000000"; 
      when 941 => DO <= x"00000000"; 
      when 942 => DO <= x"00000000"; 
      when 943 => DO <= x"00000000"; 
      when 944 => DO <= x"00000000"; 
      when 945 => DO <= x"00000000"; 
      when 946 => DO <= x"00000000"; 
      when 947 => DO <= x"00000000"; 
      when 948 => DO <= x"00000000"; 
      when 949 => DO <= x"00000000"; 
      when 950 => DO <= x"00000000"; 
      when 951 => DO <= x"00000000"; 
      when 952 => DO <= x"00000000"; 
      when 953 => DO <= x"00000000"; 
      when 954 => DO <= x"00000000"; 
      when 955 => DO <= x"00000000"; 
      when 956 => DO <= x"00000000"; 
      when 957 => DO <= x"00000000"; 
      when 958 => DO <= x"00000000"; 
      when 959 => DO <= x"00000000"; 
      when 960 => DO <= x"00000000"; 
      when 961 => DO <= x"00000000"; 
      when 962 => DO <= x"00000000"; 
      when 963 => DO <= x"00000000"; 
      when 964 => DO <= x"00000000"; 
      when 965 => DO <= x"00000000"; 
      when 966 => DO <= x"00000000"; 
      when 967 => DO <= x"00000000"; 
      when 968 => DO <= x"00000000"; 
      when 969 => DO <= x"00000000"; 
      when 970 => DO <= x"00000000"; 
      when 971 => DO <= x"00000000"; 
      when 972 => DO <= x"00000000"; 
      when 973 => DO <= x"00000000"; 
      when 974 => DO <= x"00000000"; 
      when 975 => DO <= x"00000000"; 
      when 976 => DO <= x"00000000"; 
      when 977 => DO <= x"00000000"; 
      when 978 => DO <= x"00000000"; 
      when 979 => DO <= x"00000000"; 
      when 980 => DO <= x"00000000"; 
      when 981 => DO <= x"00000000"; 
      when 982 => DO <= x"00000000"; 
      when 983 => DO <= x"00000000"; 
      when 984 => DO <= x"00000000"; 
      when 985 => DO <= x"00000000"; 
      when 986 => DO <= x"00000000"; 
      when 987 => DO <= x"00000000"; 
      when 988 => DO <= x"00000000"; 
      when 989 => DO <= x"00000000"; 
      when 990 => DO <= x"00000000"; 
      when 991 => DO <= x"00000000"; 
      when 992 => DO <= x"00000000"; 
      when 993 => DO <= x"00000000"; 
      when 994 => DO <= x"00000000"; 
      when 995 => DO <= x"00000000"; 
      when 996 => DO <= x"00000000"; 
      when 997 => DO <= x"00000000"; 
      when 998 => DO <= x"00000000"; 
      when 999 => DO <= x"00000000"; 
      when 1000 => DO <= x"00000000"; 
      when 1001 => DO <= x"00000000"; 
      when 1002 => DO <= x"00000000"; 
      when 1003 => DO <= x"00000000"; 
      when 1004 => DO <= x"00000000"; 
      when 1005 => DO <= x"00000000"; 
      when 1006 => DO <= x"00000000"; 
      when 1007 => DO <= x"00000000"; 
      when 1008 => DO <= x"00000000"; 
      when 1009 => DO <= x"00000000"; 
      when 1010 => DO <= x"00000000"; 
      when 1011 => DO <= x"00000000"; 
      when 1012 => DO <= x"00000000"; 
      when 1013 => DO <= x"00000000"; 
      when 1014 => DO <= x"00000000"; 
      when 1015 => DO <= x"00000000"; 
      when 1016 => DO <= x"00000000"; 
      when 1017 => DO <= x"00000000"; 
      when 1018 => DO <= x"00000000"; 
      when 1019 => DO <= x"00000000"; 
      when 1020 => DO <= x"00000000"; 
      when 1021 => DO <= x"00000000"; 
      when 1022 => DO <= x"00000000"; 
      when 1023 => DO <= x"00000000"; 
      when 1024 => DO <= x"00000000"; 
      when 1025 => DO <= x"00000000"; 
      when 1026 => DO <= x"00000000"; 
      when 1027 => DO <= x"00000000"; 
      when 1028 => DO <= x"00000000"; 
      when 1029 => DO <= x"00000000"; 
      when 1030 => DO <= x"00000000"; 
      when 1031 => DO <= x"00000000"; 
      when 1032 => DO <= x"00000000"; 
      when 1033 => DO <= x"00000000"; 
      when 1034 => DO <= x"00000000"; 
      when 1035 => DO <= x"00000000"; 
      when 1036 => DO <= x"00000000"; 
      when 1037 => DO <= x"00000000"; 
      when 1038 => DO <= x"00000000"; 
      when 1039 => DO <= x"00000000"; 
      when 1040 => DO <= x"00000000"; 
      when 1041 => DO <= x"00000000"; 
      when 1042 => DO <= x"00000000"; 
      when 1043 => DO <= x"00000000"; 
      when 1044 => DO <= x"00000000"; 
      when 1045 => DO <= x"00000000"; 
      when 1046 => DO <= x"00000000"; 
      when 1047 => DO <= x"00000000"; 
      when 1048 => DO <= x"00000000"; 
      when 1049 => DO <= x"00000000"; 
      when 1050 => DO <= x"00000000"; 
      when 1051 => DO <= x"00000000"; 
      when 1052 => DO <= x"00000000"; 
      when 1053 => DO <= x"00000000"; 
      when 1054 => DO <= x"00000000"; 
      when 1055 => DO <= x"00000000"; 
      when 1056 => DO <= x"00000000"; 
      when 1057 => DO <= x"00000000"; 
      when 1058 => DO <= x"00000000"; 
      when 1059 => DO <= x"00000000"; 
      when 1060 => DO <= x"00000000"; 
      when 1061 => DO <= x"00000000"; 
      when 1062 => DO <= x"00000000"; 
      when 1063 => DO <= x"00000000"; 
      when 1064 => DO <= x"00000000"; 
      when 1065 => DO <= x"00000000"; 
      when 1066 => DO <= x"00000000"; 
      when 1067 => DO <= x"00000000"; 
      when 1068 => DO <= x"00000000"; 
      when 1069 => DO <= x"00000000"; 
      when 1070 => DO <= x"00000000"; 
      when 1071 => DO <= x"00000000"; 
      when 1072 => DO <= x"00000000"; 
      when 1073 => DO <= x"00000000"; 
      when 1074 => DO <= x"00000000"; 
      when 1075 => DO <= x"00000000"; 
      when 1076 => DO <= x"00000000"; 
      when 1077 => DO <= x"00000000"; 
      when 1078 => DO <= x"00000000"; 
      when 1079 => DO <= x"00000000"; 
      when 1080 => DO <= x"00000000"; 
      when 1081 => DO <= x"00000000"; 
      when 1082 => DO <= x"00000000"; 
      when 1083 => DO <= x"00000000"; 
      when 1084 => DO <= x"00000000"; 
      when 1085 => DO <= x"00000000"; 
      when 1086 => DO <= x"00000000"; 
      when 1087 => DO <= x"00000000"; 
      when 1088 => DO <= x"00000000"; 
      when 1089 => DO <= x"00000000"; 
      when 1090 => DO <= x"00000000"; 
      when 1091 => DO <= x"00000000"; 
      when 1092 => DO <= x"00000000"; 
      when 1093 => DO <= x"00000000"; 
      when 1094 => DO <= x"00000000"; 
      when 1095 => DO <= x"00000000"; 
      when 1096 => DO <= x"00000000"; 
      when 1097 => DO <= x"00000000"; 
      when 1098 => DO <= x"00000000"; 
      when 1099 => DO <= x"00000000"; 
      when 1100 => DO <= x"00000000"; 
      when 1101 => DO <= x"00000000"; 
      when 1102 => DO <= x"00000000"; 
      when 1103 => DO <= x"00000000"; 
      when 1104 => DO <= x"00000000"; 
      when 1105 => DO <= x"00000000"; 
      when 1106 => DO <= x"00000000"; 
      when 1107 => DO <= x"00000000"; 
      when 1108 => DO <= x"00000000"; 
      when 1109 => DO <= x"00000000"; 
      when 1110 => DO <= x"00000000"; 
      when 1111 => DO <= x"00000000"; 
      when 1112 => DO <= x"00000000"; 
      when 1113 => DO <= x"00000000"; 
      when 1114 => DO <= x"00000000"; 
      when 1115 => DO <= x"00000000"; 
      when 1116 => DO <= x"00000000"; 
      when 1117 => DO <= x"00000000"; 
      when 1118 => DO <= x"00000000"; 
      when 1119 => DO <= x"00000000"; 
      when 1120 => DO <= x"00000000"; 
      when 1121 => DO <= x"00000000"; 
      when 1122 => DO <= x"00000000"; 
      when 1123 => DO <= x"00000000"; 
      when 1124 => DO <= x"00000000"; 
      when 1125 => DO <= x"00000000"; 
      when 1126 => DO <= x"00000000"; 
      when 1127 => DO <= x"00000000"; 
      when 1128 => DO <= x"00000000"; 
      when 1129 => DO <= x"00000000"; 
      when 1130 => DO <= x"00000000"; 
      when 1131 => DO <= x"00000000"; 
      when 1132 => DO <= x"00000000"; 
      when 1133 => DO <= x"00000000"; 
      when 1134 => DO <= x"00000000"; 
      when 1135 => DO <= x"00000000"; 
      when 1136 => DO <= x"00000000"; 
      when 1137 => DO <= x"00000000"; 
      when 1138 => DO <= x"00000000"; 
      when 1139 => DO <= x"00000000"; 
      when 1140 => DO <= x"00000000"; 
      when 1141 => DO <= x"00000000"; 
      when 1142 => DO <= x"00000000"; 
      when 1143 => DO <= x"00000000"; 
      when 1144 => DO <= x"00000000"; 
      when 1145 => DO <= x"00000000"; 
      when 1146 => DO <= x"00000000"; 
      when 1147 => DO <= x"00000000"; 
      when 1148 => DO <= x"00000000"; 
      when 1149 => DO <= x"00000000"; 
      when 1150 => DO <= x"00000000"; 
      when 1151 => DO <= x"00000000"; 
      when 1152 => DO <= x"00000000"; 
      when 1153 => DO <= x"00000000"; 
      when 1154 => DO <= x"00000000"; 
      when 1155 => DO <= x"00000000"; 
      when 1156 => DO <= x"00000000"; 
      when 1157 => DO <= x"00000000"; 
      when 1158 => DO <= x"00000000"; 
      when 1159 => DO <= x"00000000"; 
      when 1160 => DO <= x"00000000"; 
      when 1161 => DO <= x"00000000"; 
      when 1162 => DO <= x"00000000"; 
      when 1163 => DO <= x"00000000"; 
      when 1164 => DO <= x"00000000"; 
      when 1165 => DO <= x"00000000"; 
      when 1166 => DO <= x"00000000"; 
      when 1167 => DO <= x"00000000"; 
      when 1168 => DO <= x"00000000"; 
      when 1169 => DO <= x"00000000"; 
      when 1170 => DO <= x"00000000"; 
      when 1171 => DO <= x"00000000"; 
      when 1172 => DO <= x"00000000"; 
      when 1173 => DO <= x"00000000"; 
      when 1174 => DO <= x"00000000"; 
      when 1175 => DO <= x"00000000"; 
      when 1176 => DO <= x"00000000"; 
      when 1177 => DO <= x"00000000"; 
      when 1178 => DO <= x"00000000"; 
      when 1179 => DO <= x"00000000"; 
      when 1180 => DO <= x"00000000"; 
      when 1181 => DO <= x"00000000"; 
      when 1182 => DO <= x"00000000"; 
      when 1183 => DO <= x"00000000"; 
      when 1184 => DO <= x"00000000"; 
      when 1185 => DO <= x"00000000"; 
      when 1186 => DO <= x"00000000"; 
      when 1187 => DO <= x"00000000"; 
      when 1188 => DO <= x"00000000"; 
      when 1189 => DO <= x"00000000"; 
      when 1190 => DO <= x"00000000"; 
      when 1191 => DO <= x"00000000"; 
      when 1192 => DO <= x"00000000"; 
      when 1193 => DO <= x"00000000"; 
      when 1194 => DO <= x"00000000"; 
      when 1195 => DO <= x"00000000"; 
      when 1196 => DO <= x"00000000"; 
      when 1197 => DO <= x"00000000"; 
      when 1198 => DO <= x"00000000"; 
      when 1199 => DO <= x"00000000"; 
      when 1200 => DO <= x"00000000"; 
      when 1201 => DO <= x"00000000"; 
      when 1202 => DO <= x"00000000"; 
      when 1203 => DO <= x"00000000"; 
      when 1204 => DO <= x"00000000"; 
      when 1205 => DO <= x"00000000"; 
      when 1206 => DO <= x"00000000"; 
      when 1207 => DO <= x"00000000"; 
      when 1208 => DO <= x"00000000"; 
      when 1209 => DO <= x"00000000"; 
      when 1210 => DO <= x"00000000"; 
      when 1211 => DO <= x"00000000"; 
      when 1212 => DO <= x"00000000"; 
      when 1213 => DO <= x"00000000"; 
      when 1214 => DO <= x"00000000"; 
      when 1215 => DO <= x"00000000"; 
      when 1216 => DO <= x"00000000"; 
      when 1217 => DO <= x"00000000"; 
      when 1218 => DO <= x"00000000"; 
      when 1219 => DO <= x"00000000"; 
      when 1220 => DO <= x"00000000"; 
      when 1221 => DO <= x"00000000"; 
      when 1222 => DO <= x"00000000"; 
      when 1223 => DO <= x"00000000"; 
      when 1224 => DO <= x"00000000"; 
      when 1225 => DO <= x"00000000"; 
      when 1226 => DO <= x"00000000"; 
      when 1227 => DO <= x"00000000"; 
      when 1228 => DO <= x"00000000"; 
      when 1229 => DO <= x"00000000"; 
      when 1230 => DO <= x"00000000"; 
      when 1231 => DO <= x"00000000"; 
      when 1232 => DO <= x"00000000"; 
      when 1233 => DO <= x"00000000"; 
      when 1234 => DO <= x"00000000"; 
      when 1235 => DO <= x"00000000"; 
      when 1236 => DO <= x"00000000"; 
      when 1237 => DO <= x"00000000"; 
      when 1238 => DO <= x"00000000"; 
      when 1239 => DO <= x"00000000"; 
      when 1240 => DO <= x"00000000"; 
      when 1241 => DO <= x"00000000"; 
      when 1242 => DO <= x"00000000"; 
      when 1243 => DO <= x"00000000"; 
      when 1244 => DO <= x"00000000"; 
      when 1245 => DO <= x"00000000"; 
      when 1246 => DO <= x"00000000"; 
      when 1247 => DO <= x"00000000"; 
      when 1248 => DO <= x"00000000"; 
      when 1249 => DO <= x"00000000"; 
      when 1250 => DO <= x"00000000"; 
      when 1251 => DO <= x"00000000"; 
      when 1252 => DO <= x"00000000"; 
      when 1253 => DO <= x"00000000"; 
      when 1254 => DO <= x"00000000"; 
      when 1255 => DO <= x"00000000"; 
      when 1256 => DO <= x"00000000"; 
      when 1257 => DO <= x"00000000"; 
      when 1258 => DO <= x"00000000"; 
      when 1259 => DO <= x"00000000"; 
      when 1260 => DO <= x"00000000"; 
      when 1261 => DO <= x"00000000"; 
      when 1262 => DO <= x"00000000"; 
      when 1263 => DO <= x"00000000"; 
      when 1264 => DO <= x"00000000"; 
      when 1265 => DO <= x"00000000"; 
      when 1266 => DO <= x"00000000"; 
      when 1267 => DO <= x"00000000"; 
      when 1268 => DO <= x"00000000"; 
      when 1269 => DO <= x"00000000"; 
      when 1270 => DO <= x"00000000"; 
      when 1271 => DO <= x"00000000"; 
      when 1272 => DO <= x"00000000"; 
      when 1273 => DO <= x"00000000"; 
      when 1274 => DO <= x"00000000"; 
      when 1275 => DO <= x"00000000"; 
      when 1276 => DO <= x"00000000"; 
      when 1277 => DO <= x"00000000"; 
      when 1278 => DO <= x"00000000"; 
      when 1279 => DO <= x"00000000"; 
      when 1280 => DO <= x"00000000"; 
      when 1281 => DO <= x"00000000"; 
      when 1282 => DO <= x"00000000"; 
      when 1283 => DO <= x"00000000"; 
      when 1284 => DO <= x"00000000"; 
      when 1285 => DO <= x"00000000"; 
      when 1286 => DO <= x"00000000"; 
      when 1287 => DO <= x"00000000"; 
      when 1288 => DO <= x"00000000"; 
      when 1289 => DO <= x"00000000"; 
      when 1290 => DO <= x"00000000"; 
      when 1291 => DO <= x"00000000"; 
      when 1292 => DO <= x"00000000"; 
      when 1293 => DO <= x"00000000"; 
      when 1294 => DO <= x"00000000"; 
      when 1295 => DO <= x"00000000"; 
      when 1296 => DO <= x"00000000"; 
      when 1297 => DO <= x"00000000"; 
      when 1298 => DO <= x"00000000"; 
      when 1299 => DO <= x"00000000"; 
      when 1300 => DO <= x"00000000"; 
      when 1301 => DO <= x"00000000"; 
      when 1302 => DO <= x"00000000"; 
      when 1303 => DO <= x"00000000"; 
      when 1304 => DO <= x"00000000"; 
      when 1305 => DO <= x"00000000"; 
      when 1306 => DO <= x"00000000"; 
      when 1307 => DO <= x"00000000"; 
      when 1308 => DO <= x"00000000"; 
      when 1309 => DO <= x"00000000"; 
      when 1310 => DO <= x"00000000"; 
      when 1311 => DO <= x"00000000"; 
      when 1312 => DO <= x"00000000"; 
      when 1313 => DO <= x"00000000"; 
      when 1314 => DO <= x"00000000"; 
      when 1315 => DO <= x"00000000"; 
      when 1316 => DO <= x"00000000"; 
      when 1317 => DO <= x"00000000"; 
      when 1318 => DO <= x"00000000"; 
      when 1319 => DO <= x"00000000"; 
      when 1320 => DO <= x"00000000"; 
      when 1321 => DO <= x"00000000"; 
      when 1322 => DO <= x"00000000"; 
      when 1323 => DO <= x"00000000"; 
      when 1324 => DO <= x"00000000"; 
      when 1325 => DO <= x"00000000"; 
      when 1326 => DO <= x"00000000"; 
      when 1327 => DO <= x"00000000"; 
      when 1328 => DO <= x"00000000"; 
      when 1329 => DO <= x"00000000"; 
      when 1330 => DO <= x"00000000"; 
      when 1331 => DO <= x"00000000"; 
      when 1332 => DO <= x"00000000"; 
      when 1333 => DO <= x"00000000"; 
      when 1334 => DO <= x"00000000"; 
      when 1335 => DO <= x"00000000"; 
      when 1336 => DO <= x"00000000"; 
      when 1337 => DO <= x"00000000"; 
      when 1338 => DO <= x"00000000"; 
      when 1339 => DO <= x"00000000"; 
      when 1340 => DO <= x"00000000"; 
      when 1341 => DO <= x"00000000"; 
      when 1342 => DO <= x"00000000"; 
      when 1343 => DO <= x"00000000"; 
      when 1344 => DO <= x"00000000"; 
      when 1345 => DO <= x"00000000"; 
      when 1346 => DO <= x"00000000"; 
      when 1347 => DO <= x"00000000"; 
      when 1348 => DO <= x"00000000"; 
      when 1349 => DO <= x"00000000"; 
      when 1350 => DO <= x"00000000"; 
      when 1351 => DO <= x"00000000"; 
      when 1352 => DO <= x"00000000"; 
      when 1353 => DO <= x"00000000"; 
      when 1354 => DO <= x"00000000"; 
      when 1355 => DO <= x"00000000"; 
      when 1356 => DO <= x"00000000"; 
      when 1357 => DO <= x"00000000"; 
      when 1358 => DO <= x"00000000"; 
      when 1359 => DO <= x"00000000"; 
      when 1360 => DO <= x"00000000"; 
      when 1361 => DO <= x"00000000"; 
      when 1362 => DO <= x"00000000"; 
      when 1363 => DO <= x"00000000"; 
      when 1364 => DO <= x"00000000"; 
      when 1365 => DO <= x"00000000"; 
      when 1366 => DO <= x"00000000"; 
      when 1367 => DO <= x"00000000"; 
      when 1368 => DO <= x"00000000"; 
      when 1369 => DO <= x"00000000"; 
      when 1370 => DO <= x"00000000"; 
      when 1371 => DO <= x"00000000"; 
      when 1372 => DO <= x"00000000"; 
      when 1373 => DO <= x"00000000"; 
      when 1374 => DO <= x"00000000"; 
      when 1375 => DO <= x"00000000"; 
      when 1376 => DO <= x"00000000"; 
      when 1377 => DO <= x"00000000"; 
      when 1378 => DO <= x"00000000"; 
      when 1379 => DO <= x"00000000"; 
      when 1380 => DO <= x"00000000"; 
      when 1381 => DO <= x"00000000"; 
      when 1382 => DO <= x"00000000"; 
      when 1383 => DO <= x"00000000"; 
      when 1384 => DO <= x"00000000"; 
      when 1385 => DO <= x"00000000"; 
      when 1386 => DO <= x"00000000"; 
      when 1387 => DO <= x"00000000"; 
      when 1388 => DO <= x"00000000"; 
      when 1389 => DO <= x"00000000"; 
      when 1390 => DO <= x"00000000"; 
      when 1391 => DO <= x"00000000"; 
      when 1392 => DO <= x"00000000"; 
      when 1393 => DO <= x"00000000"; 
      when 1394 => DO <= x"00000000"; 
      when 1395 => DO <= x"00000000"; 
      when 1396 => DO <= x"00000000"; 
      when 1397 => DO <= x"00000000"; 
      when 1398 => DO <= x"00000000"; 
      when 1399 => DO <= x"00000000"; 
      when 1400 => DO <= x"00000000"; 
      when 1401 => DO <= x"00000000"; 
      when 1402 => DO <= x"00000000"; 
      when 1403 => DO <= x"00000000"; 
      when 1404 => DO <= x"00000000"; 
      when 1405 => DO <= x"00000000"; 
      when 1406 => DO <= x"00000000"; 
      when 1407 => DO <= x"00000000"; 
      when 1408 => DO <= x"00000000"; 
      when 1409 => DO <= x"00000000"; 
      when 1410 => DO <= x"00000000"; 
      when 1411 => DO <= x"00000000"; 
      when 1412 => DO <= x"00000000"; 
      when 1413 => DO <= x"00000000"; 
      when 1414 => DO <= x"00000000"; 
      when 1415 => DO <= x"00000000"; 
      when 1416 => DO <= x"00000000"; 
      when 1417 => DO <= x"00000000"; 
      when 1418 => DO <= x"00000000"; 
      when 1419 => DO <= x"00000000"; 
      when 1420 => DO <= x"00000000"; 
      when 1421 => DO <= x"00000000"; 
      when 1422 => DO <= x"00000000"; 
      when 1423 => DO <= x"00000000"; 
      when 1424 => DO <= x"00000000"; 
      when 1425 => DO <= x"00000000"; 
      when 1426 => DO <= x"00000000"; 
      when 1427 => DO <= x"00000000"; 
      when 1428 => DO <= x"00000000"; 
      when 1429 => DO <= x"00000000"; 
      when 1430 => DO <= x"00000000"; 
      when 1431 => DO <= x"00000000"; 
      when 1432 => DO <= x"00000000"; 
      when 1433 => DO <= x"00000000"; 
      when 1434 => DO <= x"00000000"; 
      when 1435 => DO <= x"00000000"; 
      when 1436 => DO <= x"00000000"; 
      when 1437 => DO <= x"00000000"; 
      when 1438 => DO <= x"00000000"; 
      when 1439 => DO <= x"00000000"; 
      when 1440 => DO <= x"00000000"; 
      when 1441 => DO <= x"00000000"; 
      when 1442 => DO <= x"00000000"; 
      when 1443 => DO <= x"00000000"; 
      when 1444 => DO <= x"00000000"; 
      when 1445 => DO <= x"00000000"; 
      when 1446 => DO <= x"00000000"; 
      when 1447 => DO <= x"00000000"; 
      when 1448 => DO <= x"00000000"; 
      when 1449 => DO <= x"00000000"; 
      when 1450 => DO <= x"00000000"; 
      when 1451 => DO <= x"00000000"; 
      when 1452 => DO <= x"00000000"; 
      when 1453 => DO <= x"00000000"; 
      when 1454 => DO <= x"00000000"; 
      when 1455 => DO <= x"00000000"; 
      when 1456 => DO <= x"00000000"; 
      when 1457 => DO <= x"00000000"; 
      when 1458 => DO <= x"00000000"; 
      when 1459 => DO <= x"00000000"; 
      when 1460 => DO <= x"00000000"; 
      when 1461 => DO <= x"00000000"; 
      when 1462 => DO <= x"00000000"; 
      when 1463 => DO <= x"00000000"; 
      when 1464 => DO <= x"00000000"; 
      when 1465 => DO <= x"00000000"; 
      when 1466 => DO <= x"00000000"; 
      when 1467 => DO <= x"00000000"; 
      when 1468 => DO <= x"00000000"; 
      when 1469 => DO <= x"00000000"; 
      when 1470 => DO <= x"00000000"; 
      when 1471 => DO <= x"00000000"; 
      when 1472 => DO <= x"00000000"; 
      when 1473 => DO <= x"00000000"; 
      when 1474 => DO <= x"00000000"; 
      when 1475 => DO <= x"00000000"; 
      when 1476 => DO <= x"00000000"; 
      when 1477 => DO <= x"00000000"; 
      when 1478 => DO <= x"00000000"; 
      when 1479 => DO <= x"00000000"; 
      when 1480 => DO <= x"00000000"; 
      when 1481 => DO <= x"00000000"; 
      when 1482 => DO <= x"00000000"; 
      when 1483 => DO <= x"00000000"; 
      when 1484 => DO <= x"00000000"; 
      when 1485 => DO <= x"00000000"; 
      when 1486 => DO <= x"00000000"; 
      when 1487 => DO <= x"00000000"; 
      when 1488 => DO <= x"00000000"; 
      when 1489 => DO <= x"00000000"; 
      when 1490 => DO <= x"00000000"; 
      when 1491 => DO <= x"00000000"; 
      when 1492 => DO <= x"00000000"; 
      when 1493 => DO <= x"00000000"; 
      when 1494 => DO <= x"00000000"; 
      when 1495 => DO <= x"00000000"; 
      when 1496 => DO <= x"00000000"; 
      when 1497 => DO <= x"00000000"; 
      when 1498 => DO <= x"00000000"; 
      when 1499 => DO <= x"00000000"; 
      when 1500 => DO <= x"00000000"; 
      when 1501 => DO <= x"00000000"; 
      when 1502 => DO <= x"00000000"; 
      when 1503 => DO <= x"00000000"; 
      when 1504 => DO <= x"00000000"; 
      when 1505 => DO <= x"00000000"; 
      when 1506 => DO <= x"00000000"; 
      when 1507 => DO <= x"00000000"; 
      when 1508 => DO <= x"00000000"; 
      when 1509 => DO <= x"00000000"; 
      when 1510 => DO <= x"00000000"; 
      when 1511 => DO <= x"00000000"; 
      when 1512 => DO <= x"00000000"; 
      when 1513 => DO <= x"00000000"; 
      when 1514 => DO <= x"00000000"; 
      when 1515 => DO <= x"00000000"; 
      when 1516 => DO <= x"00000000"; 
      when 1517 => DO <= x"00000000"; 
      when 1518 => DO <= x"00000000"; 
      when 1519 => DO <= x"00000000"; 
      when 1520 => DO <= x"00000000"; 
      when 1521 => DO <= x"00000000"; 
      when 1522 => DO <= x"00000000"; 
      when 1523 => DO <= x"00000000"; 
      when 1524 => DO <= x"00000000"; 
      when 1525 => DO <= x"00000000"; 
      when 1526 => DO <= x"00000000"; 
      when 1527 => DO <= x"00000000"; 
      when 1528 => DO <= x"00000000"; 
      when 1529 => DO <= x"00000000"; 
      when 1530 => DO <= x"00000000"; 
      when 1531 => DO <= x"00000000"; 
      when 1532 => DO <= x"00000000"; 
      when 1533 => DO <= x"00000000"; 
      when 1534 => DO <= x"00000000"; 
      when 1535 => DO <= x"00000000"; 
      when 1536 => DO <= x"00000000"; 
      when 1537 => DO <= x"00000000"; 
      when 1538 => DO <= x"00000000"; 
      when 1539 => DO <= x"00000000"; 
      when 1540 => DO <= x"00000000"; 
      when 1541 => DO <= x"00000000"; 
      when 1542 => DO <= x"00000000"; 
      when 1543 => DO <= x"00000000"; 
      when 1544 => DO <= x"00000000"; 
      when 1545 => DO <= x"00000000"; 
      when 1546 => DO <= x"00000000"; 
      when 1547 => DO <= x"00000000"; 
      when 1548 => DO <= x"00000000"; 
      when 1549 => DO <= x"00000000"; 
      when 1550 => DO <= x"00000000"; 
      when 1551 => DO <= x"00000000"; 
      when 1552 => DO <= x"00000000"; 
      when 1553 => DO <= x"00000000"; 
      when 1554 => DO <= x"00000000"; 
      when 1555 => DO <= x"00000000"; 
      when 1556 => DO <= x"00000000"; 
      when 1557 => DO <= x"00000000"; 
      when 1558 => DO <= x"00000000"; 
      when 1559 => DO <= x"00000000"; 
      when 1560 => DO <= x"00000000"; 
      when 1561 => DO <= x"00000000"; 
      when 1562 => DO <= x"00000000"; 
      when 1563 => DO <= x"00000000"; 
      when 1564 => DO <= x"00000000"; 
      when 1565 => DO <= x"00000000"; 
      when 1566 => DO <= x"00000000"; 
      when 1567 => DO <= x"00000000"; 
      when 1568 => DO <= x"00000000"; 
      when 1569 => DO <= x"00000000"; 
      when 1570 => DO <= x"00000000"; 
      when 1571 => DO <= x"00000000"; 
      when 1572 => DO <= x"00000000"; 
      when 1573 => DO <= x"00000000"; 
      when 1574 => DO <= x"00000000"; 
      when 1575 => DO <= x"00000000"; 
      when 1576 => DO <= x"00000000"; 
      when 1577 => DO <= x"00000000"; 
      when 1578 => DO <= x"00000000"; 
      when 1579 => DO <= x"00000000"; 
      when 1580 => DO <= x"00000000"; 
      when 1581 => DO <= x"00000000"; 
      when 1582 => DO <= x"00000000"; 
      when 1583 => DO <= x"00000000"; 
      when 1584 => DO <= x"00000000"; 
      when 1585 => DO <= x"00000000"; 
      when 1586 => DO <= x"00000000"; 
      when 1587 => DO <= x"00000000"; 
      when 1588 => DO <= x"00000000"; 
      when 1589 => DO <= x"00000000"; 
      when 1590 => DO <= x"00000000"; 
      when 1591 => DO <= x"00000000"; 
      when 1592 => DO <= x"00000000"; 
      when 1593 => DO <= x"00000000"; 
      when 1594 => DO <= x"00000000"; 
      when 1595 => DO <= x"00000000"; 
      when 1596 => DO <= x"00000000"; 
      when 1597 => DO <= x"00000000"; 
      when 1598 => DO <= x"00000000"; 
      when 1599 => DO <= x"00000000"; 
      when 1600 => DO <= x"00000000"; 
      when 1601 => DO <= x"00000000"; 
      when 1602 => DO <= x"00000000"; 
      when 1603 => DO <= x"00000000"; 
      when 1604 => DO <= x"00000000"; 
      when 1605 => DO <= x"00000000"; 
      when 1606 => DO <= x"00000000"; 
      when 1607 => DO <= x"00000000"; 
      when 1608 => DO <= x"00000000"; 
      when 1609 => DO <= x"00000000"; 
      when 1610 => DO <= x"00000000"; 
      when 1611 => DO <= x"00000000"; 
      when 1612 => DO <= x"00000000"; 
      when 1613 => DO <= x"00000000"; 
      when 1614 => DO <= x"00000000"; 
      when 1615 => DO <= x"00000000"; 
      when 1616 => DO <= x"00000000"; 
      when 1617 => DO <= x"00000000"; 
      when 1618 => DO <= x"00000000"; 
      when 1619 => DO <= x"00000000"; 
      when 1620 => DO <= x"00000000"; 
      when 1621 => DO <= x"00000000"; 
      when 1622 => DO <= x"00000000"; 
      when 1623 => DO <= x"00000000"; 
      when 1624 => DO <= x"00000000"; 
      when 1625 => DO <= x"00000000"; 
      when 1626 => DO <= x"00000000"; 
      when 1627 => DO <= x"00000000"; 
      when 1628 => DO <= x"00000000"; 
      when 1629 => DO <= x"00000000"; 
      when 1630 => DO <= x"00000000"; 
      when 1631 => DO <= x"00000000"; 
      when 1632 => DO <= x"00000000"; 
      when 1633 => DO <= x"00000000"; 
      when 1634 => DO <= x"00000000"; 
      when 1635 => DO <= x"00000000"; 
      when 1636 => DO <= x"00000000"; 
      when 1637 => DO <= x"00000000"; 
      when 1638 => DO <= x"00000000"; 
      when 1639 => DO <= x"00000000"; 
      when 1640 => DO <= x"00000000"; 
      when 1641 => DO <= x"00000000"; 
      when 1642 => DO <= x"00000000"; 
      when 1643 => DO <= x"00000000"; 
      when 1644 => DO <= x"00000000"; 
      when 1645 => DO <= x"00000000"; 
      when 1646 => DO <= x"00000000"; 
      when 1647 => DO <= x"00000000"; 
      when 1648 => DO <= x"00000000"; 
      when 1649 => DO <= x"00000000"; 
      when 1650 => DO <= x"00000000"; 
      when 1651 => DO <= x"00000000"; 
      when 1652 => DO <= x"00000000"; 
      when 1653 => DO <= x"00000000"; 
      when 1654 => DO <= x"00000000"; 
      when 1655 => DO <= x"00000000"; 
      when 1656 => DO <= x"00000000"; 
      when 1657 => DO <= x"00000000"; 
      when 1658 => DO <= x"00000000"; 
      when 1659 => DO <= x"00000000"; 
      when 1660 => DO <= x"00000000"; 
      when 1661 => DO <= x"00000000"; 
      when 1662 => DO <= x"00000000"; 
      when 1663 => DO <= x"00000000"; 
      when 1664 => DO <= x"00000000"; 
      when 1665 => DO <= x"00000000"; 
      when 1666 => DO <= x"00000000"; 
      when 1667 => DO <= x"00000000"; 
      when 1668 => DO <= x"00000000"; 
      when 1669 => DO <= x"00000000"; 
      when 1670 => DO <= x"00000000"; 
      when 1671 => DO <= x"00000000"; 
      when 1672 => DO <= x"00000000"; 
      when 1673 => DO <= x"00000000"; 
      when 1674 => DO <= x"00000000"; 
      when 1675 => DO <= x"00000000"; 
      when 1676 => DO <= x"00000000"; 
      when 1677 => DO <= x"00000000"; 
      when 1678 => DO <= x"00000000"; 
      when 1679 => DO <= x"00000000"; 
      when 1680 => DO <= x"00000000"; 
      when 1681 => DO <= x"00000000"; 
      when 1682 => DO <= x"00000000"; 
      when 1683 => DO <= x"00000000"; 
      when 1684 => DO <= x"00000000"; 
      when 1685 => DO <= x"00000000"; 
      when 1686 => DO <= x"00000000"; 
      when 1687 => DO <= x"00000000"; 
      when 1688 => DO <= x"00000000"; 
      when 1689 => DO <= x"00000000"; 
      when 1690 => DO <= x"00000000"; 
      when 1691 => DO <= x"00000000"; 
      when 1692 => DO <= x"00000000"; 
      when 1693 => DO <= x"00000000"; 
      when 1694 => DO <= x"00000000"; 
      when 1695 => DO <= x"00000000"; 
      when 1696 => DO <= x"00000000"; 
      when 1697 => DO <= x"00000000"; 
      when 1698 => DO <= x"00000000"; 
      when 1699 => DO <= x"00000000"; 
      when 1700 => DO <= x"00000000"; 
      when 1701 => DO <= x"00000000"; 
      when 1702 => DO <= x"00000000"; 
      when 1703 => DO <= x"00000000"; 
      when 1704 => DO <= x"00000000"; 
      when 1705 => DO <= x"00000000"; 
      when 1706 => DO <= x"00000000"; 
      when 1707 => DO <= x"00000000"; 
      when 1708 => DO <= x"00000000"; 
      when 1709 => DO <= x"00000000"; 
      when 1710 => DO <= x"00000000"; 
      when 1711 => DO <= x"00000000"; 
      when 1712 => DO <= x"00000000"; 
      when 1713 => DO <= x"00000000"; 
      when 1714 => DO <= x"00000000"; 
      when 1715 => DO <= x"00000000"; 
      when 1716 => DO <= x"00000000"; 
      when 1717 => DO <= x"00000000"; 
      when 1718 => DO <= x"00000000"; 
      when 1719 => DO <= x"00000000"; 
      when 1720 => DO <= x"00000000"; 
      when 1721 => DO <= x"00000000"; 
      when 1722 => DO <= x"00000000"; 
      when 1723 => DO <= x"00000000"; 
      when 1724 => DO <= x"00000000"; 
      when 1725 => DO <= x"00000000"; 
      when 1726 => DO <= x"00000000"; 
      when 1727 => DO <= x"00000000"; 
      when 1728 => DO <= x"00000000"; 
      when 1729 => DO <= x"00000000"; 
      when 1730 => DO <= x"00000000"; 
      when 1731 => DO <= x"00000000"; 
      when 1732 => DO <= x"00000000"; 
      when 1733 => DO <= x"00000000"; 
      when 1734 => DO <= x"00000000"; 
      when 1735 => DO <= x"00000000"; 
      when 1736 => DO <= x"00000000"; 
      when 1737 => DO <= x"00000000"; 
      when 1738 => DO <= x"00000000"; 
      when 1739 => DO <= x"00000000"; 
      when 1740 => DO <= x"00000000"; 
      when 1741 => DO <= x"00000000"; 
      when 1742 => DO <= x"00000000"; 
      when 1743 => DO <= x"00000000"; 
      when 1744 => DO <= x"00000000"; 
      when 1745 => DO <= x"00000000"; 
      when 1746 => DO <= x"00000000"; 
      when 1747 => DO <= x"00000000"; 
      when 1748 => DO <= x"00000000"; 
      when 1749 => DO <= x"00000000"; 
      when 1750 => DO <= x"00000000"; 
      when 1751 => DO <= x"00000000"; 
      when 1752 => DO <= x"00000000"; 
      when 1753 => DO <= x"00000000"; 
      when 1754 => DO <= x"00000000"; 
      when 1755 => DO <= x"00000000"; 
      when 1756 => DO <= x"00000000"; 
      when 1757 => DO <= x"00000000"; 
      when 1758 => DO <= x"00000000"; 
      when 1759 => DO <= x"00000000"; 
      when 1760 => DO <= x"00000000"; 
      when 1761 => DO <= x"00000000"; 
      when 1762 => DO <= x"00000000"; 
      when 1763 => DO <= x"00000000"; 
      when 1764 => DO <= x"00000000"; 
      when 1765 => DO <= x"00000000"; 
      when 1766 => DO <= x"00000000"; 
      when 1767 => DO <= x"00000000"; 
      when 1768 => DO <= x"00000000"; 
      when 1769 => DO <= x"00000000"; 
      when 1770 => DO <= x"00000000"; 
      when 1771 => DO <= x"00000000"; 
      when 1772 => DO <= x"00000000"; 
      when 1773 => DO <= x"00000000"; 
      when 1774 => DO <= x"00000000"; 
      when 1775 => DO <= x"00000000"; 
      when 1776 => DO <= x"00000000"; 
      when 1777 => DO <= x"00000000"; 
      when 1778 => DO <= x"00000000"; 
      when 1779 => DO <= x"00000000"; 
      when 1780 => DO <= x"00000000"; 
      when 1781 => DO <= x"00000000"; 
      when 1782 => DO <= x"00000000"; 
      when 1783 => DO <= x"00000000"; 
      when 1784 => DO <= x"00000000"; 
      when 1785 => DO <= x"00000000"; 
      when 1786 => DO <= x"00000000"; 
      when 1787 => DO <= x"00000000"; 
      when 1788 => DO <= x"00000000"; 
      when 1789 => DO <= x"00000000"; 
      when 1790 => DO <= x"00000000"; 
      when 1791 => DO <= x"00000000"; 
      when 1792 => DO <= x"00000000"; 
      when 1793 => DO <= x"00000000"; 
      when 1794 => DO <= x"00000000"; 
      when 1795 => DO <= x"00000000"; 
      when 1796 => DO <= x"00000000"; 
      when 1797 => DO <= x"00000000"; 
      when 1798 => DO <= x"00000000"; 
      when 1799 => DO <= x"00000000"; 
      when 1800 => DO <= x"00000000"; 
      when 1801 => DO <= x"00000000"; 
      when 1802 => DO <= x"00000000"; 
      when 1803 => DO <= x"00000000"; 
      when 1804 => DO <= x"00000000"; 
      when 1805 => DO <= x"00000000"; 
      when 1806 => DO <= x"00000000"; 
      when 1807 => DO <= x"00000000"; 
      when 1808 => DO <= x"00000000"; 
      when 1809 => DO <= x"00000000"; 
      when 1810 => DO <= x"00000000"; 
      when 1811 => DO <= x"00000000"; 
      when 1812 => DO <= x"00000000"; 
      when 1813 => DO <= x"00000000"; 
      when 1814 => DO <= x"00000000"; 
      when 1815 => DO <= x"00000000"; 
      when 1816 => DO <= x"00000000"; 
      when 1817 => DO <= x"00000000"; 
      when 1818 => DO <= x"00000000"; 
      when 1819 => DO <= x"00000000"; 
      when 1820 => DO <= x"00000000"; 
      when 1821 => DO <= x"00000000"; 
      when 1822 => DO <= x"00000000"; 
      when 1823 => DO <= x"00000000"; 
      when 1824 => DO <= x"00000000"; 
      when 1825 => DO <= x"00000000"; 
      when 1826 => DO <= x"00000000"; 
      when 1827 => DO <= x"00000000"; 
      when 1828 => DO <= x"00000000"; 
      when 1829 => DO <= x"00000000"; 
      when 1830 => DO <= x"00000000"; 
      when 1831 => DO <= x"00000000"; 
      when 1832 => DO <= x"00000000"; 
      when 1833 => DO <= x"00000000"; 
      when 1834 => DO <= x"00000000"; 
      when 1835 => DO <= x"00000000"; 
      when 1836 => DO <= x"00000000"; 
      when 1837 => DO <= x"00000000"; 
      when 1838 => DO <= x"00000000"; 
      when 1839 => DO <= x"00000000"; 
      when 1840 => DO <= x"00000000"; 
      when 1841 => DO <= x"00000000"; 
      when 1842 => DO <= x"00000000"; 
      when 1843 => DO <= x"00000000"; 
      when 1844 => DO <= x"00000000"; 
      when 1845 => DO <= x"00000000"; 
      when 1846 => DO <= x"00000000"; 
      when 1847 => DO <= x"00000000"; 
      when 1848 => DO <= x"00000000"; 
      when 1849 => DO <= x"00000000"; 
      when 1850 => DO <= x"00000000"; 
      when 1851 => DO <= x"00000000"; 
      when 1852 => DO <= x"00000000"; 
      when 1853 => DO <= x"00000000"; 
      when 1854 => DO <= x"00000000"; 
      when 1855 => DO <= x"00000000"; 
      when 1856 => DO <= x"00000000"; 
      when 1857 => DO <= x"00000000"; 
      when 1858 => DO <= x"00000000"; 
      when 1859 => DO <= x"00000000"; 
      when 1860 => DO <= x"00000000"; 
      when 1861 => DO <= x"00000000"; 
      when 1862 => DO <= x"00000000"; 
      when 1863 => DO <= x"00000000"; 
      when 1864 => DO <= x"00000000"; 
      when 1865 => DO <= x"00000000"; 
      when 1866 => DO <= x"00000000"; 
      when 1867 => DO <= x"00000000"; 
      when 1868 => DO <= x"00000000"; 
      when 1869 => DO <= x"00000000"; 
      when 1870 => DO <= x"00000000"; 
      when 1871 => DO <= x"00000000"; 
      when 1872 => DO <= x"00000000"; 
      when 1873 => DO <= x"00000000"; 
      when 1874 => DO <= x"00000000"; 
      when 1875 => DO <= x"00000000"; 
      when 1876 => DO <= x"00000000"; 
      when 1877 => DO <= x"00000000"; 
      when 1878 => DO <= x"00000000"; 
      when 1879 => DO <= x"00000000"; 
      when 1880 => DO <= x"00000000"; 
      when 1881 => DO <= x"00000000"; 
      when 1882 => DO <= x"00000000"; 
      when 1883 => DO <= x"00000000"; 
      when 1884 => DO <= x"00000000"; 
      when 1885 => DO <= x"00000000"; 
      when 1886 => DO <= x"00000000"; 
      when 1887 => DO <= x"00000000"; 
      when 1888 => DO <= x"00000000"; 
      when 1889 => DO <= x"00000000"; 
      when 1890 => DO <= x"00000000"; 
      when 1891 => DO <= x"00000000"; 
      when 1892 => DO <= x"00000000"; 
      when 1893 => DO <= x"00000000"; 
      when 1894 => DO <= x"00000000"; 
      when 1895 => DO <= x"00000000"; 
      when 1896 => DO <= x"00000000"; 
      when 1897 => DO <= x"00000000"; 
      when 1898 => DO <= x"00000000"; 
      when 1899 => DO <= x"00000000"; 
      when 1900 => DO <= x"00000000"; 
      when 1901 => DO <= x"00000000"; 
      when 1902 => DO <= x"00000000"; 
      when 1903 => DO <= x"00000000"; 
      when 1904 => DO <= x"00000000"; 
      when 1905 => DO <= x"00000000"; 
      when 1906 => DO <= x"00000000"; 
      when 1907 => DO <= x"00000000"; 
      when 1908 => DO <= x"00000000"; 
      when 1909 => DO <= x"00000000"; 
      when 1910 => DO <= x"00000000"; 
      when 1911 => DO <= x"00000000"; 
      when 1912 => DO <= x"00000000"; 
      when 1913 => DO <= x"00000000"; 
      when 1914 => DO <= x"00000000"; 
      when 1915 => DO <= x"00000000"; 
      when 1916 => DO <= x"00000000"; 
      when 1917 => DO <= x"00000000"; 
      when 1918 => DO <= x"00000000"; 
      when 1919 => DO <= x"00000000"; 
      when 1920 => DO <= x"00000000"; 
      when 1921 => DO <= x"00000000"; 
      when 1922 => DO <= x"00000000"; 
      when 1923 => DO <= x"00000000"; 
      when 1924 => DO <= x"00000000"; 
      when 1925 => DO <= x"00000000"; 
      when 1926 => DO <= x"00000000"; 
      when 1927 => DO <= x"00000000"; 
      when 1928 => DO <= x"00000000"; 
      when 1929 => DO <= x"00000000"; 
      when 1930 => DO <= x"00000000"; 
      when 1931 => DO <= x"00000000"; 
      when 1932 => DO <= x"00000000"; 
      when 1933 => DO <= x"00000000"; 
      when 1934 => DO <= x"00000000"; 
      when 1935 => DO <= x"00000000"; 
      when 1936 => DO <= x"00000000"; 
      when 1937 => DO <= x"00000000"; 
      when 1938 => DO <= x"00000000"; 
      when 1939 => DO <= x"00000000"; 
      when 1940 => DO <= x"00000000"; 
      when 1941 => DO <= x"00000000"; 
      when 1942 => DO <= x"00000000"; 
      when 1943 => DO <= x"00000000"; 
      when 1944 => DO <= x"00000000"; 
      when 1945 => DO <= x"00000000"; 
      when 1946 => DO <= x"00000000"; 
      when 1947 => DO <= x"00000000"; 
      when 1948 => DO <= x"00000000"; 
      when 1949 => DO <= x"00000000"; 
      when 1950 => DO <= x"00000000"; 
      when 1951 => DO <= x"00000000"; 
      when 1952 => DO <= x"00000000"; 
      when 1953 => DO <= x"00000000"; 
      when 1954 => DO <= x"00000000"; 
      when 1955 => DO <= x"00000000"; 
      when 1956 => DO <= x"00000000"; 
      when 1957 => DO <= x"00000000"; 
      when 1958 => DO <= x"00000000"; 
      when 1959 => DO <= x"00000000"; 
      when 1960 => DO <= x"00000000"; 
      when 1961 => DO <= x"00000000"; 
      when 1962 => DO <= x"00000000"; 
      when 1963 => DO <= x"00000000"; 
      when 1964 => DO <= x"00000000"; 
      when 1965 => DO <= x"00000000"; 
      when 1966 => DO <= x"00000000"; 
      when 1967 => DO <= x"00000000"; 
      when 1968 => DO <= x"00000000"; 
      when 1969 => DO <= x"00000000"; 
      when 1970 => DO <= x"00000000"; 
      when 1971 => DO <= x"00000000"; 
      when 1972 => DO <= x"00000000"; 
      when 1973 => DO <= x"00000000"; 
      when 1974 => DO <= x"00000000"; 
      when 1975 => DO <= x"00000000"; 
      when 1976 => DO <= x"00000000"; 
      when 1977 => DO <= x"00000000"; 
      when 1978 => DO <= x"00000000"; 
      when 1979 => DO <= x"00000000"; 
      when 1980 => DO <= x"00000000"; 
      when 1981 => DO <= x"00000000"; 
      when 1982 => DO <= x"00000000"; 
      when 1983 => DO <= x"00000000"; 
      when 1984 => DO <= x"00000000"; 
      when 1985 => DO <= x"00000000"; 
      when 1986 => DO <= x"00000000"; 
      when 1987 => DO <= x"00000000"; 
      when 1988 => DO <= x"00000000"; 
      when 1989 => DO <= x"00000000"; 
      when 1990 => DO <= x"00000000"; 
      when 1991 => DO <= x"00000000"; 
      when 1992 => DO <= x"00000000"; 
      when 1993 => DO <= x"00000000"; 
      when 1994 => DO <= x"00000000"; 
      when 1995 => DO <= x"00000000"; 
      when 1996 => DO <= x"00000000"; 
      when 1997 => DO <= x"00000000"; 
      when 1998 => DO <= x"00000000"; 
      when 1999 => DO <= x"00000000"; 
      when 2000 => DO <= x"00000000"; 
      when 2001 => DO <= x"00000000"; 
      when 2002 => DO <= x"00000000"; 
      when 2003 => DO <= x"00000000"; 
      when 2004 => DO <= x"00000000"; 
      when 2005 => DO <= x"00000000"; 
      when 2006 => DO <= x"00000000"; 
      when 2007 => DO <= x"00000000"; 
      when 2008 => DO <= x"00000000"; 
      when 2009 => DO <= x"00000000"; 
      when 2010 => DO <= x"00000000"; 
      when 2011 => DO <= x"00000000"; 
      when 2012 => DO <= x"00000000"; 
      when 2013 => DO <= x"00000000"; 
      when 2014 => DO <= x"00000000"; 
      when 2015 => DO <= x"00000000"; 
      when 2016 => DO <= x"00000000"; 
      when 2017 => DO <= x"00000000"; 
      when 2018 => DO <= x"00000000"; 
      when 2019 => DO <= x"00000000"; 
      when 2020 => DO <= x"00000000"; 
      when 2021 => DO <= x"00000000"; 
      when 2022 => DO <= x"00000000"; 
      when 2023 => DO <= x"00000000"; 
      when 2024 => DO <= x"00000000"; 
      when 2025 => DO <= x"00000000"; 
      when 2026 => DO <= x"00000000"; 
      when 2027 => DO <= x"00000000"; 
      when 2028 => DO <= x"00000000"; 
      when 2029 => DO <= x"00000000"; 
      when 2030 => DO <= x"00000000"; 
      when 2031 => DO <= x"00000000"; 
      when 2032 => DO <= x"00000000"; 
      when 2033 => DO <= x"00000000"; 
      when 2034 => DO <= x"00000000"; 
      when 2035 => DO <= x"00000000"; 
      when 2036 => DO <= x"00000000"; 
      when 2037 => DO <= x"00000000"; 
      when 2038 => DO <= x"00000000"; 
      when 2039 => DO <= x"00000000"; 
      when 2040 => DO <= x"00000000"; 
      when 2041 => DO <= x"00000000"; 
      when 2042 => DO <= x"00000000"; 
      when 2043 => DO <= x"00000000"; 
      when 2044 => DO <= x"00000000"; 
      when 2045 => DO <= x"00000000"; 
      when 2046 => DO <= x"00000000"; 
      when 2047 => DO <= x"00000000"; 
      when 2048 => DO <= x"00000000"; 
      when 2049 => DO <= x"00000000"; 
      when 2050 => DO <= x"00000000"; 
      when 2051 => DO <= x"00000000"; 
      when 2052 => DO <= x"00000000"; 
      when 2053 => DO <= x"00000000"; 
      when 2054 => DO <= x"00000000"; 
      when 2055 => DO <= x"00000000"; 
      when 2056 => DO <= x"00000000"; 
      when 2057 => DO <= x"00000000"; 
      when 2058 => DO <= x"00000000"; 
      when 2059 => DO <= x"00000000"; 
      when 2060 => DO <= x"00000000"; 
      when 2061 => DO <= x"00000000"; 
      when 2062 => DO <= x"00000000"; 
      when 2063 => DO <= x"00000000"; 
      when 2064 => DO <= x"00000000"; 
      when 2065 => DO <= x"00000000"; 
      when 2066 => DO <= x"00000000"; 
      when 2067 => DO <= x"00000000"; 
      when 2068 => DO <= x"00000000"; 
      when 2069 => DO <= x"00000000"; 
      when 2070 => DO <= x"00000000"; 
      when 2071 => DO <= x"00000000"; 
      when 2072 => DO <= x"00000000"; 
      when 2073 => DO <= x"00000000"; 
      when 2074 => DO <= x"00000000"; 
      when 2075 => DO <= x"00000000"; 
      when 2076 => DO <= x"00000000"; 
      when 2077 => DO <= x"00000000"; 
      when 2078 => DO <= x"00000000"; 
      when 2079 => DO <= x"00000000"; 
      when 2080 => DO <= x"00000000"; 
      when 2081 => DO <= x"00000000"; 
      when 2082 => DO <= x"00000000"; 
      when 2083 => DO <= x"00000000"; 
      when 2084 => DO <= x"00000000"; 
      when 2085 => DO <= x"00000000"; 
      when 2086 => DO <= x"00000000"; 
      when 2087 => DO <= x"00000000"; 
      when 2088 => DO <= x"00000000"; 
      when 2089 => DO <= x"00000000"; 
      when 2090 => DO <= x"00000000"; 
      when 2091 => DO <= x"00000000"; 
      when 2092 => DO <= x"00000000"; 
      when 2093 => DO <= x"00000000"; 
      when 2094 => DO <= x"00000000"; 
      when 2095 => DO <= x"00000000"; 
      when 2096 => DO <= x"00000000"; 
      when 2097 => DO <= x"00000000"; 
      when 2098 => DO <= x"00000000"; 
      when 2099 => DO <= x"00000000"; 
      when 2100 => DO <= x"00000000"; 
      when 2101 => DO <= x"00000000"; 
      when 2102 => DO <= x"00000000"; 
      when 2103 => DO <= x"00000000"; 
      when 2104 => DO <= x"00000000"; 
      when 2105 => DO <= x"00000000"; 
      when 2106 => DO <= x"00000000"; 
      when 2107 => DO <= x"00000000"; 
      when 2108 => DO <= x"00000000"; 
      when 2109 => DO <= x"00000000"; 
      when 2110 => DO <= x"00000000"; 
      when 2111 => DO <= x"00000000"; 
      when 2112 => DO <= x"00000000"; 
      when 2113 => DO <= x"00000000"; 
      when 2114 => DO <= x"00000000"; 
      when 2115 => DO <= x"00000000"; 
      when 2116 => DO <= x"00000000"; 
      when 2117 => DO <= x"00000000"; 
      when 2118 => DO <= x"00000000"; 
      when 2119 => DO <= x"00000000"; 
      when 2120 => DO <= x"00000000"; 
      when 2121 => DO <= x"00000000"; 
      when 2122 => DO <= x"00000000"; 
      when 2123 => DO <= x"00000000"; 
      when 2124 => DO <= x"00000000"; 
      when 2125 => DO <= x"00000000"; 
      when 2126 => DO <= x"00000000"; 
      when 2127 => DO <= x"00000000"; 
      when 2128 => DO <= x"00000000"; 
      when 2129 => DO <= x"00000000"; 
      when 2130 => DO <= x"00000000"; 
      when 2131 => DO <= x"00000000"; 
      when 2132 => DO <= x"00000000"; 
      when 2133 => DO <= x"00000000"; 
      when 2134 => DO <= x"00000000"; 
      when 2135 => DO <= x"00000000"; 
      when 2136 => DO <= x"00000000"; 
      when 2137 => DO <= x"00000000"; 
      when 2138 => DO <= x"00000000"; 
      when 2139 => DO <= x"00000000"; 
      when 2140 => DO <= x"00000000"; 
      when 2141 => DO <= x"00000000"; 
      when 2142 => DO <= x"00000000"; 
      when 2143 => DO <= x"00000000"; 
      when 2144 => DO <= x"00000000"; 
      when 2145 => DO <= x"00000000"; 
      when 2146 => DO <= x"00000000"; 
      when 2147 => DO <= x"00000000"; 
      when 2148 => DO <= x"00000000"; 
      when 2149 => DO <= x"00000000"; 
      when 2150 => DO <= x"00000000"; 
      when 2151 => DO <= x"00000000"; 
      when 2152 => DO <= x"00000000"; 
      when 2153 => DO <= x"00000000"; 
      when 2154 => DO <= x"00000000"; 
      when 2155 => DO <= x"00000000"; 
      when 2156 => DO <= x"00000000"; 
      when 2157 => DO <= x"00000000"; 
      when 2158 => DO <= x"00000000"; 
      when 2159 => DO <= x"00000000"; 
      when 2160 => DO <= x"00000000"; 
      when 2161 => DO <= x"00000000"; 
      when 2162 => DO <= x"00000000"; 
      when 2163 => DO <= x"00000000"; 
      when 2164 => DO <= x"00000000"; 
      when 2165 => DO <= x"00000000"; 
      when 2166 => DO <= x"00000000"; 
      when 2167 => DO <= x"00000000"; 
      when 2168 => DO <= x"00000000"; 
      when 2169 => DO <= x"00000000"; 
      when 2170 => DO <= x"00000000"; 
      when 2171 => DO <= x"00000000"; 
      when 2172 => DO <= x"00000000"; 
      when 2173 => DO <= x"00000000"; 
      when 2174 => DO <= x"00000000"; 
      when 2175 => DO <= x"00000000"; 
      when 2176 => DO <= x"00000000"; 
      when 2177 => DO <= x"00000000"; 
      when 2178 => DO <= x"00000000"; 
      when 2179 => DO <= x"00000000"; 
      when 2180 => DO <= x"00000000"; 
      when 2181 => DO <= x"00000000"; 
      when 2182 => DO <= x"00000000"; 
      when 2183 => DO <= x"00000000"; 
      when 2184 => DO <= x"00000000"; 
      when 2185 => DO <= x"00000000"; 
      when 2186 => DO <= x"00000000"; 
      when 2187 => DO <= x"00000000"; 
      when 2188 => DO <= x"00000000"; 
      when 2189 => DO <= x"00000000"; 
      when 2190 => DO <= x"00000000"; 
      when 2191 => DO <= x"00000000"; 
      when 2192 => DO <= x"00000000"; 
      when 2193 => DO <= x"00000000"; 
      when 2194 => DO <= x"00000000"; 
      when 2195 => DO <= x"00000000"; 
      when 2196 => DO <= x"00000000"; 
      when 2197 => DO <= x"00000000"; 
      when 2198 => DO <= x"00000000"; 
      when 2199 => DO <= x"00000000"; 
      when 2200 => DO <= x"00000000"; 
      when 2201 => DO <= x"00000000"; 
      when 2202 => DO <= x"00000000"; 
      when 2203 => DO <= x"00000000"; 
      when 2204 => DO <= x"00000000"; 
      when 2205 => DO <= x"00000000"; 
      when 2206 => DO <= x"00000000"; 
      when 2207 => DO <= x"00000000"; 
      when 2208 => DO <= x"00000000"; 
      when 2209 => DO <= x"00000000"; 
      when 2210 => DO <= x"00000000"; 
      when 2211 => DO <= x"00000000"; 
      when 2212 => DO <= x"00000000"; 
      when 2213 => DO <= x"00000000"; 
      when 2214 => DO <= x"00000000"; 
      when 2215 => DO <= x"00000000"; 
      when 2216 => DO <= x"00000000"; 
      when 2217 => DO <= x"00000000"; 
      when 2218 => DO <= x"00000000"; 
      when 2219 => DO <= x"00000000"; 
      when 2220 => DO <= x"00000000"; 
      when 2221 => DO <= x"00000000"; 
      when 2222 => DO <= x"00000000"; 
      when 2223 => DO <= x"00000000"; 
      when 2224 => DO <= x"00000000"; 
      when 2225 => DO <= x"00000000"; 
      when 2226 => DO <= x"00000000"; 
      when 2227 => DO <= x"00000000"; 
      when 2228 => DO <= x"00000000"; 
      when 2229 => DO <= x"00000000"; 
      when 2230 => DO <= x"00000000"; 
      when 2231 => DO <= x"00000000"; 
      when 2232 => DO <= x"00000000"; 
      when 2233 => DO <= x"00000000"; 
      when 2234 => DO <= x"00000000"; 
      when 2235 => DO <= x"00000000"; 
      when 2236 => DO <= x"00000000"; 
      when 2237 => DO <= x"00000000"; 
      when 2238 => DO <= x"00000000"; 
      when 2239 => DO <= x"00000000"; 
      when 2240 => DO <= x"00000000"; 
      when 2241 => DO <= x"00000000"; 
      when 2242 => DO <= x"00000000"; 
      when 2243 => DO <= x"00000000"; 
      when 2244 => DO <= x"00000000"; 
      when 2245 => DO <= x"00000000"; 
      when 2246 => DO <= x"00000000"; 
      when 2247 => DO <= x"00000000"; 
      when 2248 => DO <= x"00000000"; 
      when 2249 => DO <= x"00000000"; 
      when 2250 => DO <= x"00000000"; 
      when 2251 => DO <= x"00000000"; 
      when 2252 => DO <= x"00000000"; 
      when 2253 => DO <= x"00000000"; 
      when 2254 => DO <= x"00000000"; 
      when 2255 => DO <= x"00000000"; 
      when 2256 => DO <= x"00000000"; 
      when 2257 => DO <= x"00000000"; 
      when 2258 => DO <= x"00000000"; 
      when 2259 => DO <= x"00000000"; 
      when 2260 => DO <= x"00000000"; 
      when 2261 => DO <= x"00000000"; 
      when 2262 => DO <= x"00000000"; 
      when 2263 => DO <= x"00000000"; 
      when 2264 => DO <= x"00000000"; 
      when 2265 => DO <= x"00000000"; 
      when 2266 => DO <= x"00000000"; 
      when 2267 => DO <= x"00000000"; 
      when 2268 => DO <= x"00000000"; 
      when 2269 => DO <= x"00000000"; 
      when 2270 => DO <= x"00000000"; 
      when 2271 => DO <= x"00000000"; 
      when 2272 => DO <= x"00000000"; 
      when 2273 => DO <= x"00000000"; 
      when 2274 => DO <= x"00000000"; 
      when 2275 => DO <= x"00000000"; 
      when 2276 => DO <= x"00000000"; 
      when 2277 => DO <= x"00000000"; 
      when 2278 => DO <= x"00000000"; 
      when 2279 => DO <= x"00000000"; 
      when 2280 => DO <= x"00000000"; 
      when 2281 => DO <= x"00000000"; 
      when 2282 => DO <= x"00000000"; 
      when 2283 => DO <= x"00000000"; 
      when 2284 => DO <= x"00000000"; 
      when 2285 => DO <= x"00000000"; 
      when 2286 => DO <= x"00000000"; 
      when 2287 => DO <= x"00000000"; 
      when 2288 => DO <= x"00000000"; 
      when 2289 => DO <= x"00000000"; 
      when 2290 => DO <= x"00000000"; 
      when 2291 => DO <= x"00000000"; 
      when 2292 => DO <= x"00000000"; 
      when 2293 => DO <= x"00000000"; 
      when 2294 => DO <= x"00000000"; 
      when 2295 => DO <= x"00000000"; 
      when 2296 => DO <= x"00000000"; 
      when 2297 => DO <= x"00000000"; 
      when 2298 => DO <= x"00000000"; 
      when 2299 => DO <= x"00000000"; 
      when 2300 => DO <= x"00000000"; 
      when 2301 => DO <= x"00000000"; 
      when 2302 => DO <= x"00000000"; 
      when 2303 => DO <= x"00000000"; 
      when 2304 => DO <= x"00000000"; 
      when 2305 => DO <= x"00000000"; 
      when 2306 => DO <= x"00000000"; 
      when 2307 => DO <= x"00000000"; 
      when 2308 => DO <= x"00000000"; 
      when 2309 => DO <= x"00000000"; 
      when 2310 => DO <= x"00000000"; 
      when 2311 => DO <= x"00000000"; 
      when 2312 => DO <= x"00000000"; 
      when 2313 => DO <= x"00000000"; 
      when 2314 => DO <= x"00000000"; 
      when 2315 => DO <= x"00000000"; 
      when 2316 => DO <= x"00000000"; 
      when 2317 => DO <= x"00000000"; 
      when 2318 => DO <= x"00000000"; 
      when 2319 => DO <= x"00000000"; 
      when 2320 => DO <= x"00000000"; 
      when 2321 => DO <= x"00000000"; 
      when 2322 => DO <= x"00000000"; 
      when 2323 => DO <= x"00000000"; 
      when 2324 => DO <= x"00000000"; 
      when 2325 => DO <= x"00000000"; 
      when 2326 => DO <= x"00000000"; 
      when 2327 => DO <= x"00000000"; 
      when 2328 => DO <= x"00000000"; 
      when 2329 => DO <= x"00000000"; 
      when 2330 => DO <= x"00000000"; 
      when 2331 => DO <= x"00000000"; 
      when 2332 => DO <= x"00000000"; 
      when 2333 => DO <= x"00000000"; 
      when 2334 => DO <= x"00000000"; 
      when 2335 => DO <= x"00000000"; 
      when 2336 => DO <= x"00000000"; 
      when 2337 => DO <= x"00000000"; 
      when 2338 => DO <= x"00000000"; 
      when 2339 => DO <= x"00000000"; 
      when 2340 => DO <= x"00000000"; 
      when 2341 => DO <= x"00000000"; 
      when 2342 => DO <= x"00000000"; 
      when 2343 => DO <= x"00000000"; 
      when 2344 => DO <= x"00000000"; 
      when 2345 => DO <= x"00000000"; 
      when 2346 => DO <= x"00000000"; 
      when 2347 => DO <= x"00000000"; 
      when 2348 => DO <= x"00000000"; 
      when 2349 => DO <= x"00000000"; 
      when 2350 => DO <= x"00000000"; 
      when 2351 => DO <= x"00000000"; 
      when 2352 => DO <= x"00000000"; 
      when 2353 => DO <= x"00000000"; 
      when 2354 => DO <= x"00000000"; 
      when 2355 => DO <= x"00000000"; 
      when 2356 => DO <= x"00000000"; 
      when 2357 => DO <= x"00000000"; 
      when 2358 => DO <= x"00000000"; 
      when 2359 => DO <= x"00000000"; 
      when 2360 => DO <= x"00000000"; 
      when 2361 => DO <= x"00000000"; 
      when 2362 => DO <= x"00000000"; 
      when 2363 => DO <= x"00000000"; 
      when 2364 => DO <= x"00000000"; 
      when 2365 => DO <= x"00000000"; 
      when 2366 => DO <= x"00000000"; 
      when 2367 => DO <= x"00000000"; 
      when 2368 => DO <= x"00000000"; 
      when 2369 => DO <= x"00000000"; 
      when 2370 => DO <= x"00000000"; 
      when 2371 => DO <= x"00000000"; 
      when 2372 => DO <= x"00000000"; 
      when 2373 => DO <= x"00000000"; 
      when 2374 => DO <= x"00000000"; 
      when 2375 => DO <= x"00000000"; 
      when 2376 => DO <= x"00000000"; 
      when 2377 => DO <= x"00000000"; 
      when 2378 => DO <= x"00000000"; 
      when 2379 => DO <= x"00000000"; 
      when 2380 => DO <= x"00000000"; 
      when 2381 => DO <= x"00000000"; 
      when 2382 => DO <= x"00000000"; 
      when 2383 => DO <= x"00000000"; 
      when 2384 => DO <= x"00000000"; 
      when 2385 => DO <= x"00000000"; 
      when 2386 => DO <= x"00000000"; 
      when 2387 => DO <= x"00000000"; 
      when 2388 => DO <= x"00000000"; 
      when 2389 => DO <= x"00000000"; 
      when 2390 => DO <= x"00000000"; 
      when 2391 => DO <= x"00000000"; 
      when 2392 => DO <= x"00000000"; 
      when 2393 => DO <= x"00000000"; 
      when 2394 => DO <= x"00000000"; 
      when 2395 => DO <= x"00000000"; 
      when 2396 => DO <= x"00000000"; 
      when 2397 => DO <= x"00000000"; 
      when 2398 => DO <= x"00000000"; 
      when 2399 => DO <= x"00000000"; 
      when 2400 => DO <= x"00000000"; 
      when 2401 => DO <= x"00000000"; 
      when 2402 => DO <= x"00000000"; 
      when 2403 => DO <= x"00000000"; 
      when 2404 => DO <= x"00000000"; 
      when 2405 => DO <= x"00000000"; 
      when 2406 => DO <= x"00000000"; 
      when 2407 => DO <= x"00000000"; 
      when 2408 => DO <= x"00000000"; 
      when 2409 => DO <= x"00000000"; 
      when 2410 => DO <= x"00000000"; 
      when 2411 => DO <= x"00000000"; 
      when 2412 => DO <= x"00000000"; 
      when 2413 => DO <= x"00000000"; 
      when 2414 => DO <= x"00000000"; 
      when 2415 => DO <= x"00000000"; 
      when 2416 => DO <= x"00000000"; 
      when 2417 => DO <= x"00000000"; 
      when 2418 => DO <= x"00000000"; 
      when 2419 => DO <= x"00000000"; 
      when 2420 => DO <= x"00000000"; 
      when 2421 => DO <= x"00000000"; 
      when 2422 => DO <= x"00000000"; 
      when 2423 => DO <= x"00000000"; 
      when 2424 => DO <= x"00000000"; 
      when 2425 => DO <= x"00000000"; 
      when 2426 => DO <= x"00000000"; 
      when 2427 => DO <= x"00000000"; 
      when 2428 => DO <= x"00000000"; 
      when 2429 => DO <= x"00000000"; 
      when 2430 => DO <= x"00000000"; 
      when 2431 => DO <= x"00000000"; 
      when 2432 => DO <= x"00000000"; 
      when 2433 => DO <= x"00000000"; 
      when 2434 => DO <= x"00000000"; 
      when 2435 => DO <= x"00000000"; 
      when 2436 => DO <= x"00000000"; 
      when 2437 => DO <= x"00000000"; 
      when 2438 => DO <= x"00000000"; 
      when 2439 => DO <= x"00000000"; 
      when 2440 => DO <= x"00000000"; 
      when 2441 => DO <= x"00000000"; 
      when 2442 => DO <= x"00000000"; 
      when 2443 => DO <= x"00000000"; 
      when 2444 => DO <= x"00000000"; 
      when 2445 => DO <= x"00000000"; 
      when 2446 => DO <= x"00000000"; 
      when 2447 => DO <= x"00000000"; 
      when 2448 => DO <= x"00000000"; 
      when 2449 => DO <= x"00000000"; 
      when 2450 => DO <= x"00000000"; 
      when 2451 => DO <= x"00000000"; 
      when 2452 => DO <= x"00000000"; 
      when 2453 => DO <= x"00000000"; 
      when 2454 => DO <= x"00000000"; 
      when 2455 => DO <= x"00000000"; 
      when 2456 => DO <= x"00000000"; 
      when 2457 => DO <= x"00000000"; 
      when 2458 => DO <= x"00000000"; 
      when 2459 => DO <= x"00000000"; 
      when 2460 => DO <= x"00000000"; 
      when 2461 => DO <= x"00000000"; 
      when 2462 => DO <= x"00000000"; 
      when 2463 => DO <= x"00000000"; 
      when 2464 => DO <= x"00000000"; 
      when 2465 => DO <= x"00000000"; 
      when 2466 => DO <= x"00000000"; 
      when 2467 => DO <= x"00000000"; 
      when 2468 => DO <= x"00000000"; 
      when 2469 => DO <= x"00000000"; 
      when 2470 => DO <= x"00000000"; 
      when 2471 => DO <= x"00000000"; 
      when 2472 => DO <= x"00000000"; 
      when 2473 => DO <= x"00000000"; 
      when 2474 => DO <= x"00000000"; 
      when 2475 => DO <= x"00000000"; 
      when 2476 => DO <= x"00000000"; 
      when 2477 => DO <= x"00000000"; 
      when 2478 => DO <= x"00000000"; 
      when 2479 => DO <= x"00000000"; 
      when 2480 => DO <= x"00000000"; 
      when 2481 => DO <= x"00000000"; 
      when 2482 => DO <= x"00000000"; 
      when 2483 => DO <= x"00000000"; 
      when 2484 => DO <= x"00000000"; 
      when 2485 => DO <= x"00000000"; 
      when 2486 => DO <= x"00000000"; 
      when 2487 => DO <= x"00000000"; 
      when 2488 => DO <= x"00000000"; 
      when 2489 => DO <= x"00000000"; 
      when 2490 => DO <= x"00000000"; 
      when 2491 => DO <= x"00000000"; 
      when 2492 => DO <= x"00000000"; 
      when 2493 => DO <= x"00000000"; 
      when 2494 => DO <= x"00000000"; 
      when 2495 => DO <= x"00000000"; 
      when 2496 => DO <= x"00000000"; 
      when 2497 => DO <= x"00000000"; 
      when 2498 => DO <= x"00000000"; 
      when 2499 => DO <= x"00000000"; 
      when 2500 => DO <= x"00000000"; 
      when 2501 => DO <= x"00000000"; 
      when 2502 => DO <= x"00000000"; 
      when 2503 => DO <= x"00000000"; 
      when 2504 => DO <= x"00000000"; 
      when 2505 => DO <= x"00000000"; 
      when 2506 => DO <= x"00000000"; 
      when 2507 => DO <= x"00000000"; 
      when 2508 => DO <= x"00000000"; 
      when 2509 => DO <= x"00000000"; 
      when 2510 => DO <= x"00000000"; 
      when 2511 => DO <= x"00000000"; 
      when 2512 => DO <= x"00000000"; 
      when 2513 => DO <= x"00000000"; 
      when 2514 => DO <= x"00000000"; 
      when 2515 => DO <= x"00000000"; 
      when 2516 => DO <= x"00000000"; 
      when 2517 => DO <= x"00000000"; 
      when 2518 => DO <= x"00000000"; 
      when 2519 => DO <= x"00000000"; 
      when 2520 => DO <= x"00000000"; 
      when 2521 => DO <= x"00000000"; 
      when 2522 => DO <= x"00000000"; 
      when 2523 => DO <= x"00000000"; 
      when 2524 => DO <= x"00000000"; 
      when 2525 => DO <= x"00000000"; 
      when 2526 => DO <= x"00000000"; 
      when 2527 => DO <= x"00000000"; 
      when 2528 => DO <= x"00000000"; 
      when 2529 => DO <= x"00000000"; 
      when 2530 => DO <= x"00000000"; 
      when 2531 => DO <= x"00000000"; 
      when 2532 => DO <= x"00000000"; 
      when 2533 => DO <= x"00000000"; 
      when 2534 => DO <= x"00000000"; 
      when 2535 => DO <= x"00000000"; 
      when 2536 => DO <= x"00000000"; 
      when 2537 => DO <= x"00000000"; 
      when 2538 => DO <= x"00000000"; 
      when 2539 => DO <= x"00000000"; 
      when 2540 => DO <= x"00000000"; 
      when 2541 => DO <= x"00000000"; 
      when 2542 => DO <= x"00000000"; 
      when 2543 => DO <= x"00000000"; 
      when 2544 => DO <= x"00000000"; 
      when 2545 => DO <= x"00000000"; 
      when 2546 => DO <= x"00000000"; 
      when 2547 => DO <= x"00000000"; 
      when 2548 => DO <= x"00000000"; 
      when 2549 => DO <= x"00000000"; 
      when 2550 => DO <= x"00000000"; 
      when 2551 => DO <= x"00000000"; 
      when 2552 => DO <= x"00000000"; 
      when 2553 => DO <= x"00000000"; 
      when 2554 => DO <= x"00000000"; 
      when 2555 => DO <= x"00000000"; 
      when 2556 => DO <= x"00000000"; 
      when 2557 => DO <= x"00000000"; 
      when 2558 => DO <= x"00000000"; 
      when 2559 => DO <= x"00000000"; 
      when 2560 => DO <= x"00000000"; 
      when 2561 => DO <= x"00000000"; 
      when 2562 => DO <= x"00000000"; 
      when 2563 => DO <= x"00000000"; 
      when 2564 => DO <= x"00000000"; 
      when 2565 => DO <= x"00000000"; 
      when 2566 => DO <= x"00000000"; 
      when 2567 => DO <= x"00000000"; 
      when 2568 => DO <= x"00000000"; 
      when 2569 => DO <= x"00000000"; 
      when 2570 => DO <= x"00000000"; 
      when 2571 => DO <= x"00000000"; 
      when 2572 => DO <= x"00000000"; 
      when 2573 => DO <= x"00000000"; 
      when 2574 => DO <= x"00000000"; 
      when 2575 => DO <= x"00000000"; 
      when 2576 => DO <= x"00000000"; 
      when 2577 => DO <= x"00000000"; 
      when 2578 => DO <= x"00000000"; 
      when 2579 => DO <= x"00000000"; 
      when 2580 => DO <= x"00000000"; 
      when 2581 => DO <= x"00000000"; 
      when 2582 => DO <= x"00000000"; 
      when 2583 => DO <= x"00000000"; 
      when 2584 => DO <= x"00000000"; 
      when 2585 => DO <= x"00000000"; 
      when 2586 => DO <= x"00000000"; 
      when 2587 => DO <= x"00000000"; 
      when 2588 => DO <= x"00000000"; 
      when 2589 => DO <= x"00000000"; 
      when 2590 => DO <= x"00000000"; 
      when 2591 => DO <= x"00000000"; 
      when 2592 => DO <= x"00000000"; 
      when 2593 => DO <= x"00000000"; 
      when 2594 => DO <= x"00000000"; 
      when 2595 => DO <= x"00000000"; 
      when 2596 => DO <= x"00000000"; 
      when 2597 => DO <= x"00000000"; 
      when 2598 => DO <= x"00000000"; 
      when 2599 => DO <= x"00000000"; 
      when 2600 => DO <= x"00000000"; 
      when 2601 => DO <= x"00000000"; 
      when 2602 => DO <= x"00000000"; 
      when 2603 => DO <= x"00000000"; 
      when 2604 => DO <= x"00000000"; 
      when 2605 => DO <= x"00000000"; 
      when 2606 => DO <= x"00000000"; 
      when 2607 => DO <= x"00000000"; 
      when 2608 => DO <= x"00000000"; 
      when 2609 => DO <= x"00000000"; 
      when 2610 => DO <= x"00000000"; 
      when 2611 => DO <= x"00000000"; 
      when 2612 => DO <= x"00000000"; 
      when 2613 => DO <= x"00000000"; 
      when 2614 => DO <= x"00000000"; 
      when 2615 => DO <= x"00000000"; 
      when 2616 => DO <= x"00000000"; 
      when 2617 => DO <= x"00000000"; 
      when 2618 => DO <= x"00000000"; 
      when 2619 => DO <= x"00000000"; 
      when 2620 => DO <= x"00000000"; 
      when 2621 => DO <= x"00000000"; 
      when 2622 => DO <= x"00000000"; 
      when 2623 => DO <= x"00000000"; 
      when 2624 => DO <= x"00000000"; 
      when 2625 => DO <= x"00000000"; 
      when 2626 => DO <= x"00000000"; 
      when 2627 => DO <= x"00000000"; 
      when 2628 => DO <= x"00000000"; 
      when 2629 => DO <= x"00000000"; 
      when 2630 => DO <= x"00000000"; 
      when 2631 => DO <= x"00000000"; 
      when 2632 => DO <= x"00000000"; 
      when 2633 => DO <= x"00000000"; 
      when 2634 => DO <= x"00000000"; 
      when 2635 => DO <= x"00000000"; 
      when 2636 => DO <= x"00000000"; 
      when 2637 => DO <= x"00000000"; 
      when 2638 => DO <= x"00000000"; 
      when 2639 => DO <= x"00000000"; 
      when 2640 => DO <= x"00000000"; 
      when 2641 => DO <= x"00000000"; 
      when 2642 => DO <= x"00000000"; 
      when 2643 => DO <= x"00000000"; 
      when 2644 => DO <= x"00000000"; 
      when 2645 => DO <= x"00000000"; 
      when 2646 => DO <= x"00000000"; 
      when 2647 => DO <= x"00000000"; 
      when 2648 => DO <= x"00000000"; 
      when 2649 => DO <= x"00000000"; 
      when 2650 => DO <= x"00000000"; 
      when 2651 => DO <= x"00000000"; 
      when 2652 => DO <= x"00000000"; 
      when 2653 => DO <= x"00000000"; 
      when 2654 => DO <= x"00000000"; 
      when 2655 => DO <= x"00000000"; 
      when 2656 => DO <= x"00000000"; 
      when 2657 => DO <= x"00000000"; 
      when 2658 => DO <= x"00000000"; 
      when 2659 => DO <= x"00000000"; 
      when 2660 => DO <= x"00000000"; 
      when 2661 => DO <= x"00000000"; 
      when 2662 => DO <= x"00000000"; 
      when 2663 => DO <= x"00000000"; 
      when 2664 => DO <= x"00000000"; 
      when 2665 => DO <= x"00000000"; 
      when 2666 => DO <= x"00000000"; 
      when 2667 => DO <= x"00000000"; 
      when 2668 => DO <= x"00000000"; 
      when 2669 => DO <= x"00000000"; 
      when 2670 => DO <= x"00000000"; 
      when 2671 => DO <= x"00000000"; 
      when 2672 => DO <= x"00000000"; 
      when 2673 => DO <= x"00000000"; 
      when 2674 => DO <= x"00000000"; 
      when 2675 => DO <= x"00000000"; 
      when 2676 => DO <= x"00000000"; 
      when 2677 => DO <= x"00000000"; 
      when 2678 => DO <= x"00000000"; 
      when 2679 => DO <= x"00000000"; 
      when 2680 => DO <= x"00000000"; 
      when 2681 => DO <= x"00000000"; 
      when 2682 => DO <= x"00000000"; 
      when 2683 => DO <= x"00000000"; 
      when 2684 => DO <= x"00000000"; 
      when 2685 => DO <= x"00000000"; 
      when 2686 => DO <= x"00000000"; 
      when 2687 => DO <= x"00000000"; 
      when 2688 => DO <= x"00000000"; 
      when 2689 => DO <= x"00000000"; 
      when 2690 => DO <= x"00000000"; 
      when 2691 => DO <= x"00000000"; 
      when 2692 => DO <= x"00000000"; 
      when 2693 => DO <= x"00000000"; 
      when 2694 => DO <= x"00000000"; 
      when 2695 => DO <= x"00000000"; 
      when 2696 => DO <= x"00000000"; 
      when 2697 => DO <= x"00000000"; 
      when 2698 => DO <= x"00000000"; 
      when 2699 => DO <= x"00000000"; 
      when 2700 => DO <= x"00000000"; 
      when 2701 => DO <= x"00000000"; 
      when 2702 => DO <= x"00000000"; 
      when 2703 => DO <= x"00000000"; 
      when 2704 => DO <= x"00000000"; 
      when 2705 => DO <= x"00000000"; 
      when 2706 => DO <= x"00000000"; 
      when 2707 => DO <= x"00000000"; 
      when 2708 => DO <= x"00000000"; 
      when 2709 => DO <= x"00000000"; 
      when 2710 => DO <= x"00000000"; 
      when 2711 => DO <= x"00000000"; 
      when 2712 => DO <= x"00000000"; 
      when 2713 => DO <= x"00000000"; 
      when 2714 => DO <= x"00000000"; 
      when 2715 => DO <= x"00000000"; 
      when 2716 => DO <= x"00000000"; 
      when 2717 => DO <= x"00000000"; 
      when 2718 => DO <= x"00000000"; 
      when 2719 => DO <= x"00000000"; 
      when 2720 => DO <= x"00000000"; 
      when 2721 => DO <= x"00000000"; 
      when 2722 => DO <= x"00000000"; 
      when 2723 => DO <= x"00000000"; 
      when 2724 => DO <= x"00000000"; 
      when 2725 => DO <= x"00000000"; 
      when 2726 => DO <= x"00000000"; 
      when 2727 => DO <= x"00000000"; 
      when 2728 => DO <= x"00000000"; 
      when 2729 => DO <= x"00000000"; 
      when 2730 => DO <= x"00000000"; 
      when 2731 => DO <= x"00000000"; 
      when 2732 => DO <= x"00000000"; 
      when 2733 => DO <= x"00000000"; 
      when 2734 => DO <= x"00000000"; 
      when 2735 => DO <= x"00000000"; 
      when 2736 => DO <= x"00000000"; 
      when 2737 => DO <= x"00000000"; 
      when 2738 => DO <= x"00000000"; 
      when 2739 => DO <= x"00000000"; 
      when 2740 => DO <= x"00000000"; 
      when 2741 => DO <= x"00000000"; 
      when 2742 => DO <= x"00000000"; 
      when 2743 => DO <= x"00000000"; 
      when 2744 => DO <= x"00000000"; 
      when 2745 => DO <= x"00000000"; 
      when 2746 => DO <= x"00000000"; 
      when 2747 => DO <= x"00000000"; 
      when 2748 => DO <= x"00000000"; 
      when 2749 => DO <= x"00000000"; 
      when 2750 => DO <= x"00000000"; 
      when 2751 => DO <= x"00000000"; 
      when 2752 => DO <= x"00000000"; 
      when 2753 => DO <= x"00000000"; 
      when 2754 => DO <= x"00000000"; 
      when 2755 => DO <= x"00000000"; 
      when 2756 => DO <= x"00000000"; 
      when 2757 => DO <= x"00000000"; 
      when 2758 => DO <= x"00000000"; 
      when 2759 => DO <= x"00000000"; 
      when 2760 => DO <= x"00000000"; 
      when 2761 => DO <= x"00000000"; 
      when 2762 => DO <= x"00000000"; 
      when 2763 => DO <= x"00000000"; 
      when 2764 => DO <= x"00000000"; 
      when 2765 => DO <= x"00000000"; 
      when 2766 => DO <= x"00000000"; 
      when 2767 => DO <= x"00000000"; 
      when 2768 => DO <= x"00000000"; 
      when 2769 => DO <= x"00000000"; 
      when 2770 => DO <= x"00000000"; 
      when 2771 => DO <= x"00000000"; 
      when 2772 => DO <= x"00000000"; 
      when 2773 => DO <= x"00000000"; 
      when 2774 => DO <= x"00000000"; 
      when 2775 => DO <= x"00000000"; 
      when 2776 => DO <= x"00000000"; 
      when 2777 => DO <= x"00000000"; 
      when 2778 => DO <= x"00000000"; 
      when 2779 => DO <= x"00000000"; 
      when 2780 => DO <= x"00000000"; 
      when 2781 => DO <= x"00000000"; 
      when 2782 => DO <= x"00000000"; 
      when 2783 => DO <= x"00000000"; 
      when 2784 => DO <= x"00000000"; 
      when 2785 => DO <= x"00000000"; 
      when 2786 => DO <= x"00000000"; 
      when 2787 => DO <= x"00000000"; 
      when 2788 => DO <= x"00000000"; 
      when 2789 => DO <= x"00000000"; 
      when 2790 => DO <= x"00000000"; 
      when 2791 => DO <= x"00000000"; 
      when 2792 => DO <= x"00000000"; 
      when 2793 => DO <= x"00000000"; 
      when 2794 => DO <= x"00000000"; 
      when 2795 => DO <= x"00000000"; 
      when 2796 => DO <= x"00000000"; 
      when 2797 => DO <= x"00000000"; 
      when 2798 => DO <= x"00000000"; 
      when 2799 => DO <= x"00000000"; 
      when 2800 => DO <= x"00000000"; 
      when 2801 => DO <= x"00000000"; 
      when 2802 => DO <= x"00000000"; 
      when 2803 => DO <= x"00000000"; 
      when 2804 => DO <= x"00000000"; 
      when 2805 => DO <= x"00000000"; 
      when 2806 => DO <= x"00000000"; 
      when 2807 => DO <= x"00000000"; 
      when 2808 => DO <= x"00000000"; 
      when 2809 => DO <= x"00000000"; 
      when 2810 => DO <= x"00000000"; 
      when 2811 => DO <= x"00000000"; 
      when 2812 => DO <= x"00000000"; 
      when 2813 => DO <= x"00000000"; 
      when 2814 => DO <= x"00000000"; 
      when 2815 => DO <= x"00000000"; 
      when 2816 => DO <= x"00000000"; 
      when 2817 => DO <= x"00000000"; 
      when 2818 => DO <= x"00000000"; 
      when 2819 => DO <= x"00000000"; 
      when 2820 => DO <= x"00000000"; 
      when 2821 => DO <= x"00000000"; 
      when 2822 => DO <= x"00000000"; 
      when 2823 => DO <= x"00000000"; 
      when 2824 => DO <= x"00000000"; 
      when 2825 => DO <= x"00000000"; 
      when 2826 => DO <= x"00000000"; 
      when 2827 => DO <= x"00000000"; 
      when 2828 => DO <= x"00000000"; 
      when 2829 => DO <= x"00000000"; 
      when 2830 => DO <= x"00000000"; 
      when 2831 => DO <= x"00000000"; 
      when 2832 => DO <= x"00000000"; 
      when 2833 => DO <= x"00000000"; 
      when 2834 => DO <= x"00000000"; 
      when 2835 => DO <= x"00000000"; 
      when 2836 => DO <= x"00000000"; 
      when 2837 => DO <= x"00000000"; 
      when 2838 => DO <= x"00000000"; 
      when 2839 => DO <= x"00000000"; 
      when 2840 => DO <= x"00000000"; 
      when 2841 => DO <= x"00000000"; 
      when 2842 => DO <= x"00000000"; 
      when 2843 => DO <= x"00000000"; 
      when 2844 => DO <= x"00000000"; 
      when 2845 => DO <= x"00000000"; 
      when 2846 => DO <= x"00000000"; 
      when 2847 => DO <= x"00000000"; 
      when 2848 => DO <= x"00000000"; 
      when 2849 => DO <= x"00000000"; 
      when 2850 => DO <= x"00000000"; 
      when 2851 => DO <= x"00000000"; 
      when 2852 => DO <= x"00000000"; 
      when 2853 => DO <= x"00000000"; 
      when 2854 => DO <= x"00000000"; 
      when 2855 => DO <= x"00000000"; 
      when 2856 => DO <= x"00000000"; 
      when 2857 => DO <= x"00000000"; 
      when 2858 => DO <= x"00000000"; 
      when 2859 => DO <= x"00000000"; 
      when 2860 => DO <= x"00000000"; 
      when 2861 => DO <= x"00000000"; 
      when 2862 => DO <= x"00000000"; 
      when 2863 => DO <= x"00000000"; 
      when 2864 => DO <= x"00000000"; 
      when 2865 => DO <= x"00000000"; 
      when 2866 => DO <= x"00000000"; 
      when 2867 => DO <= x"00000000"; 
      when 2868 => DO <= x"00000000"; 
      when 2869 => DO <= x"00000000"; 
      when 2870 => DO <= x"00000000"; 
      when 2871 => DO <= x"00000000"; 
      when 2872 => DO <= x"00000000"; 
      when 2873 => DO <= x"00000000"; 
      when 2874 => DO <= x"00000000"; 
      when 2875 => DO <= x"00000000"; 
      when 2876 => DO <= x"00000000"; 
      when 2877 => DO <= x"00000000"; 
      when 2878 => DO <= x"00000000"; 
      when 2879 => DO <= x"00000000"; 
      when 2880 => DO <= x"00000000"; 
      when 2881 => DO <= x"00000000"; 
      when 2882 => DO <= x"00000000"; 
      when 2883 => DO <= x"00000000"; 
      when 2884 => DO <= x"00000000"; 
      when 2885 => DO <= x"00000000"; 
      when 2886 => DO <= x"00000000"; 
      when 2887 => DO <= x"00000000"; 
      when 2888 => DO <= x"00000000"; 
      when 2889 => DO <= x"00000000"; 
      when 2890 => DO <= x"00000000"; 
      when 2891 => DO <= x"00000000"; 
      when 2892 => DO <= x"00000000"; 
      when 2893 => DO <= x"00000000"; 
      when 2894 => DO <= x"00000000"; 
      when 2895 => DO <= x"00000000"; 
      when 2896 => DO <= x"00000000"; 
      when 2897 => DO <= x"00000000"; 
      when 2898 => DO <= x"00000000"; 
      when 2899 => DO <= x"00000000"; 
      when 2900 => DO <= x"00000000"; 
      when 2901 => DO <= x"00000000"; 
      when 2902 => DO <= x"00000000"; 
      when 2903 => DO <= x"00000000"; 
      when 2904 => DO <= x"00000000"; 
      when 2905 => DO <= x"00000000"; 
      when 2906 => DO <= x"00000000"; 
      when 2907 => DO <= x"00000000"; 
      when 2908 => DO <= x"00000000"; 
      when 2909 => DO <= x"00000000"; 
      when 2910 => DO <= x"00000000"; 
      when 2911 => DO <= x"00000000"; 
      when 2912 => DO <= x"00000000"; 
      when 2913 => DO <= x"00000000"; 
      when 2914 => DO <= x"00000000"; 
      when 2915 => DO <= x"00000000"; 
      when 2916 => DO <= x"00000000"; 
      when 2917 => DO <= x"00000000"; 
      when 2918 => DO <= x"00000000"; 
      when 2919 => DO <= x"00000000"; 
      when 2920 => DO <= x"00000000"; 
      when 2921 => DO <= x"00000000"; 
      when 2922 => DO <= x"00000000"; 
      when 2923 => DO <= x"00000000"; 
      when 2924 => DO <= x"00000000"; 
      when 2925 => DO <= x"00000000"; 
      when 2926 => DO <= x"00000000"; 
      when 2927 => DO <= x"00000000"; 
      when 2928 => DO <= x"00000000"; 
      when 2929 => DO <= x"00000000"; 
      when 2930 => DO <= x"00000000"; 
      when 2931 => DO <= x"00000000"; 
      when 2932 => DO <= x"00000000"; 
      when 2933 => DO <= x"00000000"; 
      when 2934 => DO <= x"00000000"; 
      when 2935 => DO <= x"00000000"; 
      when 2936 => DO <= x"00000000"; 
      when 2937 => DO <= x"00000000"; 
      when 2938 => DO <= x"00000000"; 
      when 2939 => DO <= x"00000000"; 
      when 2940 => DO <= x"00000000"; 
      when 2941 => DO <= x"00000000"; 
      when 2942 => DO <= x"00000000"; 
      when 2943 => DO <= x"00000000"; 
      when 2944 => DO <= x"00000000"; 
      when 2945 => DO <= x"00000000"; 
      when 2946 => DO <= x"00000000"; 
      when 2947 => DO <= x"00000000"; 
      when 2948 => DO <= x"00000000"; 
      when 2949 => DO <= x"00000000"; 
      when 2950 => DO <= x"00000000"; 
      when 2951 => DO <= x"00000000"; 
      when 2952 => DO <= x"00000000"; 
      when 2953 => DO <= x"00000000"; 
      when 2954 => DO <= x"00000000"; 
      when 2955 => DO <= x"00000000"; 
      when 2956 => DO <= x"00000000"; 
      when 2957 => DO <= x"00000000"; 
      when 2958 => DO <= x"00000000"; 
      when 2959 => DO <= x"00000000"; 
      when 2960 => DO <= x"00000000"; 
      when 2961 => DO <= x"00000000"; 
      when 2962 => DO <= x"00000000"; 
      when 2963 => DO <= x"00000000"; 
      when 2964 => DO <= x"00000000"; 
      when 2965 => DO <= x"00000000"; 
      when 2966 => DO <= x"00000000"; 
      when 2967 => DO <= x"00000000"; 
      when 2968 => DO <= x"00000000"; 
      when 2969 => DO <= x"00000000"; 
      when 2970 => DO <= x"00000000"; 
      when 2971 => DO <= x"00000000"; 
      when 2972 => DO <= x"00000000"; 
      when 2973 => DO <= x"00000000"; 
      when 2974 => DO <= x"00000000"; 
      when 2975 => DO <= x"00000000"; 
      when 2976 => DO <= x"00000000"; 
      when 2977 => DO <= x"00000000"; 
      when 2978 => DO <= x"00000000"; 
      when 2979 => DO <= x"00000000"; 
      when 2980 => DO <= x"00000000"; 
      when 2981 => DO <= x"00000000"; 
      when 2982 => DO <= x"00000000"; 
      when 2983 => DO <= x"00000000"; 
      when 2984 => DO <= x"00000000"; 
      when 2985 => DO <= x"00000000"; 
      when 2986 => DO <= x"00000000"; 
      when 2987 => DO <= x"00000000"; 
      when 2988 => DO <= x"00000000"; 
      when 2989 => DO <= x"00000000"; 
      when 2990 => DO <= x"00000000"; 
      when 2991 => DO <= x"00000000"; 
      when 2992 => DO <= x"00000000"; 
      when 2993 => DO <= x"00000000"; 
      when 2994 => DO <= x"00000000"; 
      when 2995 => DO <= x"00000000"; 
      when 2996 => DO <= x"00000000"; 
      when 2997 => DO <= x"00000000"; 
      when 2998 => DO <= x"00000000"; 
      when 2999 => DO <= x"00000000"; 
      when 3000 => DO <= x"00000000"; 
      when 3001 => DO <= x"00000000"; 
      when 3002 => DO <= x"00000000"; 
      when 3003 => DO <= x"00000000"; 
      when 3004 => DO <= x"00000000"; 
      when 3005 => DO <= x"00000000"; 
      when 3006 => DO <= x"00000000"; 
      when 3007 => DO <= x"00000000"; 
      when 3008 => DO <= x"00000000"; 
      when 3009 => DO <= x"00000000"; 
      when 3010 => DO <= x"00000000"; 
      when 3011 => DO <= x"00000000"; 
      when 3012 => DO <= x"00000000"; 
      when 3013 => DO <= x"00000000"; 
      when 3014 => DO <= x"00000000"; 
      when 3015 => DO <= x"00000000"; 
      when 3016 => DO <= x"00000000"; 
      when 3017 => DO <= x"00000000"; 
      when 3018 => DO <= x"00000000"; 
      when 3019 => DO <= x"00000000"; 
      when 3020 => DO <= x"00000000"; 
      when 3021 => DO <= x"00000000"; 
      when 3022 => DO <= x"00000000"; 
      when 3023 => DO <= x"00000000"; 
      when 3024 => DO <= x"00000000"; 
      when 3025 => DO <= x"00000000"; 
      when 3026 => DO <= x"00000000"; 
      when 3027 => DO <= x"00000000"; 
      when 3028 => DO <= x"00000000"; 
      when 3029 => DO <= x"00000000"; 
      when 3030 => DO <= x"00000000"; 
      when 3031 => DO <= x"00000000"; 
      when 3032 => DO <= x"00000000"; 
      when 3033 => DO <= x"00000000"; 
      when 3034 => DO <= x"00000000"; 
      when 3035 => DO <= x"00000000"; 
      when 3036 => DO <= x"00000000"; 
      when 3037 => DO <= x"00000000"; 
      when 3038 => DO <= x"00000000"; 
      when 3039 => DO <= x"00000000"; 
      when 3040 => DO <= x"00000000"; 
      when 3041 => DO <= x"00000000"; 
      when 3042 => DO <= x"00000000"; 
      when 3043 => DO <= x"00000000"; 
      when 3044 => DO <= x"00000000"; 
      when 3045 => DO <= x"00000000"; 
      when 3046 => DO <= x"00000000"; 
      when 3047 => DO <= x"00000000"; 
      when 3048 => DO <= x"00000000"; 
      when 3049 => DO <= x"00000000"; 
      when 3050 => DO <= x"00000000"; 
      when 3051 => DO <= x"00000000"; 
      when 3052 => DO <= x"00000000"; 
      when 3053 => DO <= x"00000000"; 
      when 3054 => DO <= x"00000000"; 
      when 3055 => DO <= x"00000000"; 
      when 3056 => DO <= x"00000000"; 
      when 3057 => DO <= x"00000000"; 
      when 3058 => DO <= x"00000000"; 
      when 3059 => DO <= x"00000000"; 
      when 3060 => DO <= x"00000000"; 
      when 3061 => DO <= x"00000000"; 
      when 3062 => DO <= x"00000000"; 
      when 3063 => DO <= x"00000000"; 
      when 3064 => DO <= x"00000000"; 
      when 3065 => DO <= x"00000000"; 
      when 3066 => DO <= x"00000000"; 
      when 3067 => DO <= x"00000000"; 
      when 3068 => DO <= x"00000000"; 
      when 3069 => DO <= x"00000000"; 
      when 3070 => DO <= x"00000000"; 
      when 3071 => DO <= x"00000000"; 
      when 3072 => DO <= x"00000000"; 
      when 3073 => DO <= x"00000000"; 
      when 3074 => DO <= x"00000000"; 
      when 3075 => DO <= x"00000000"; 
      when 3076 => DO <= x"00000000"; 
      when 3077 => DO <= x"00000000"; 
      when 3078 => DO <= x"00000000"; 
      when 3079 => DO <= x"00000000"; 
      when 3080 => DO <= x"00000000"; 
      when 3081 => DO <= x"00000000"; 
      when 3082 => DO <= x"00000000"; 
      when 3083 => DO <= x"00000000"; 
      when 3084 => DO <= x"00000000"; 
      when 3085 => DO <= x"00000000"; 
      when 3086 => DO <= x"00000000"; 
      when 3087 => DO <= x"00000000"; 
      when 3088 => DO <= x"00000000"; 
      when 3089 => DO <= x"00000000"; 
      when 3090 => DO <= x"00000000"; 
      when 3091 => DO <= x"00000000"; 
      when 3092 => DO <= x"00000000"; 
      when 3093 => DO <= x"00000000"; 
      when 3094 => DO <= x"00000000"; 
      when 3095 => DO <= x"00000000"; 
      when 3096 => DO <= x"00000000"; 
      when 3097 => DO <= x"00000000"; 
      when 3098 => DO <= x"00000000"; 
      when 3099 => DO <= x"00000000"; 
      when 3100 => DO <= x"00000000"; 
      when 3101 => DO <= x"00000000"; 
      when 3102 => DO <= x"00000000"; 
      when 3103 => DO <= x"00000000"; 
      when 3104 => DO <= x"00000000"; 
      when 3105 => DO <= x"00000000"; 
      when 3106 => DO <= x"00000000"; 
      when 3107 => DO <= x"00000000"; 
      when 3108 => DO <= x"00000000"; 
      when 3109 => DO <= x"00000000"; 
      when 3110 => DO <= x"00000000"; 
      when 3111 => DO <= x"00000000"; 
      when 3112 => DO <= x"00000000"; 
      when 3113 => DO <= x"00000000"; 
      when 3114 => DO <= x"00000000"; 
      when 3115 => DO <= x"00000000"; 
      when 3116 => DO <= x"00000000"; 
      when 3117 => DO <= x"00000000"; 
      when 3118 => DO <= x"00000000"; 
      when 3119 => DO <= x"00000000"; 
      when 3120 => DO <= x"00000000"; 
      when 3121 => DO <= x"00000000"; 
      when 3122 => DO <= x"00000000"; 
      when 3123 => DO <= x"00000000"; 
      when 3124 => DO <= x"00000000"; 
      when 3125 => DO <= x"00000000"; 
      when 3126 => DO <= x"00000000"; 
      when 3127 => DO <= x"00000000"; 
      when 3128 => DO <= x"00000000"; 
      when 3129 => DO <= x"00000000"; 
      when 3130 => DO <= x"00000000"; 
      when 3131 => DO <= x"00000000"; 
      when 3132 => DO <= x"00000000"; 
      when 3133 => DO <= x"00000000"; 
      when 3134 => DO <= x"00000000"; 
      when 3135 => DO <= x"00000000"; 
      when 3136 => DO <= x"00000000"; 
      when 3137 => DO <= x"00000000"; 
      when 3138 => DO <= x"00000000"; 
      when 3139 => DO <= x"00000000"; 
      when 3140 => DO <= x"00000000"; 
      when 3141 => DO <= x"00000000"; 
      when 3142 => DO <= x"00000000"; 
      when 3143 => DO <= x"00000000"; 
      when 3144 => DO <= x"00000000"; 
      when 3145 => DO <= x"00000000"; 
      when 3146 => DO <= x"00000000"; 
      when 3147 => DO <= x"00000000"; 
      when 3148 => DO <= x"00000000"; 
      when 3149 => DO <= x"00000000"; 
      when 3150 => DO <= x"00000000"; 
      when 3151 => DO <= x"00000000"; 
      when 3152 => DO <= x"00000000"; 
      when 3153 => DO <= x"00000000"; 
      when 3154 => DO <= x"00000000"; 
      when 3155 => DO <= x"00000000"; 
      when 3156 => DO <= x"00000000"; 
      when 3157 => DO <= x"00000000"; 
      when 3158 => DO <= x"00000000"; 
      when 3159 => DO <= x"00000000"; 
      when 3160 => DO <= x"00000000"; 
      when 3161 => DO <= x"00000000"; 
      when 3162 => DO <= x"00000000"; 
      when 3163 => DO <= x"00000000"; 
      when 3164 => DO <= x"00000000"; 
      when 3165 => DO <= x"00000000"; 
      when 3166 => DO <= x"00000000"; 
      when 3167 => DO <= x"00000000"; 
      when 3168 => DO <= x"00000000"; 
      when 3169 => DO <= x"00000000"; 
      when 3170 => DO <= x"00000000"; 
      when 3171 => DO <= x"00000000"; 
      when 3172 => DO <= x"00000000"; 
      when 3173 => DO <= x"00000000"; 
      when 3174 => DO <= x"00000000"; 
      when 3175 => DO <= x"00000000"; 
      when 3176 => DO <= x"00000000"; 
      when 3177 => DO <= x"00000000"; 
      when 3178 => DO <= x"00000000"; 
      when 3179 => DO <= x"00000000"; 
      when 3180 => DO <= x"00000000"; 
      when 3181 => DO <= x"00000000"; 
      when 3182 => DO <= x"00000000"; 
      when 3183 => DO <= x"00000000"; 
      when 3184 => DO <= x"00000000"; 
      when 3185 => DO <= x"00000000"; 
      when 3186 => DO <= x"00000000"; 
      when 3187 => DO <= x"00000000"; 
      when 3188 => DO <= x"00000000"; 
      when 3189 => DO <= x"00000000"; 
      when 3190 => DO <= x"00000000"; 
      when 3191 => DO <= x"00000000"; 
      when 3192 => DO <= x"00000000"; 
      when 3193 => DO <= x"00000000"; 
      when 3194 => DO <= x"00000000"; 
      when 3195 => DO <= x"00000000"; 
      when 3196 => DO <= x"00000000"; 
      when 3197 => DO <= x"00000000"; 
      when 3198 => DO <= x"00000000"; 
      when 3199 => DO <= x"00000000"; 
      when 3200 => DO <= x"00000000"; 
      when 3201 => DO <= x"00000000"; 
      when 3202 => DO <= x"00000000"; 
      when 3203 => DO <= x"00000000"; 
      when 3204 => DO <= x"00000000"; 
      when 3205 => DO <= x"00000000"; 
      when 3206 => DO <= x"00000000"; 
      when 3207 => DO <= x"00000000"; 
      when 3208 => DO <= x"00000000"; 
      when 3209 => DO <= x"00000000"; 
      when 3210 => DO <= x"00000000"; 
      when 3211 => DO <= x"00000000"; 
      when 3212 => DO <= x"00000000"; 
      when 3213 => DO <= x"00000000"; 
      when 3214 => DO <= x"00000000"; 
      when 3215 => DO <= x"00000000"; 
      when 3216 => DO <= x"00000000"; 
      when 3217 => DO <= x"00000000"; 
      when 3218 => DO <= x"00000000"; 
      when 3219 => DO <= x"00000000"; 
      when 3220 => DO <= x"00000000"; 
      when 3221 => DO <= x"00000000"; 
      when 3222 => DO <= x"00000000"; 
      when 3223 => DO <= x"00000000"; 
      when 3224 => DO <= x"00000000"; 
      when 3225 => DO <= x"00000000"; 
      when 3226 => DO <= x"00000000"; 
      when 3227 => DO <= x"00000000"; 
      when 3228 => DO <= x"00000000"; 
      when 3229 => DO <= x"00000000"; 
      when 3230 => DO <= x"00000000"; 
      when 3231 => DO <= x"00000000"; 
      when 3232 => DO <= x"00000000"; 
      when 3233 => DO <= x"00000000"; 
      when 3234 => DO <= x"00000000"; 
      when 3235 => DO <= x"00000000"; 
      when 3236 => DO <= x"00000000"; 
      when 3237 => DO <= x"00000000"; 
      when 3238 => DO <= x"00000000"; 
      when 3239 => DO <= x"00000000"; 
      when 3240 => DO <= x"00000000"; 
      when 3241 => DO <= x"00000000"; 
      when 3242 => DO <= x"00000000"; 
      when 3243 => DO <= x"00000000"; 
      when 3244 => DO <= x"00000000"; 
      when 3245 => DO <= x"00000000"; 
      when 3246 => DO <= x"00000000"; 
      when 3247 => DO <= x"00000000"; 
      when 3248 => DO <= x"00000000"; 
      when 3249 => DO <= x"00000000"; 
      when 3250 => DO <= x"00000000"; 
      when 3251 => DO <= x"00000000"; 
      when 3252 => DO <= x"00000000"; 
      when 3253 => DO <= x"00000000"; 
      when 3254 => DO <= x"00000000"; 
      when 3255 => DO <= x"00000000"; 
      when 3256 => DO <= x"00000000"; 
      when 3257 => DO <= x"00000000"; 
      when 3258 => DO <= x"00000000"; 
      when 3259 => DO <= x"00000000"; 
      when 3260 => DO <= x"00000000"; 
      when 3261 => DO <= x"00000000"; 
      when 3262 => DO <= x"00000000"; 
      when 3263 => DO <= x"00000000"; 
      when 3264 => DO <= x"00000000"; 
      when 3265 => DO <= x"00000000"; 
      when 3266 => DO <= x"00000000"; 
      when 3267 => DO <= x"00000000"; 
      when 3268 => DO <= x"00000000"; 
      when 3269 => DO <= x"00000000"; 
      when 3270 => DO <= x"00000000"; 
      when 3271 => DO <= x"00000000"; 
      when 3272 => DO <= x"00000000"; 
      when 3273 => DO <= x"00000000"; 
      when 3274 => DO <= x"00000000"; 
      when 3275 => DO <= x"00000000"; 
      when 3276 => DO <= x"00000000"; 
      when 3277 => DO <= x"00000000"; 
      when 3278 => DO <= x"00000000"; 
      when 3279 => DO <= x"00000000"; 
      when 3280 => DO <= x"00000000"; 
      when 3281 => DO <= x"00000000"; 
      when 3282 => DO <= x"00000000"; 
      when 3283 => DO <= x"00000000"; 
      when 3284 => DO <= x"00000000"; 
      when 3285 => DO <= x"00000000"; 
      when 3286 => DO <= x"00000000"; 
      when 3287 => DO <= x"00000000"; 
      when 3288 => DO <= x"00000000"; 
      when 3289 => DO <= x"00000000"; 
      when 3290 => DO <= x"00000000"; 
      when 3291 => DO <= x"00000000"; 
      when 3292 => DO <= x"00000000"; 
      when 3293 => DO <= x"00000000"; 
      when 3294 => DO <= x"00000000"; 
      when 3295 => DO <= x"00000000"; 
      when 3296 => DO <= x"00000000"; 
      when 3297 => DO <= x"00000000"; 
      when 3298 => DO <= x"00000000"; 
      when 3299 => DO <= x"00000000"; 
      when 3300 => DO <= x"00000000"; 
      when 3301 => DO <= x"00000000"; 
      when 3302 => DO <= x"00000000"; 
      when 3303 => DO <= x"00000000"; 
      when 3304 => DO <= x"00000000"; 
      when 3305 => DO <= x"00000000"; 
      when 3306 => DO <= x"00000000"; 
      when 3307 => DO <= x"00000000"; 
      when 3308 => DO <= x"00000000"; 
      when 3309 => DO <= x"00000000"; 
      when 3310 => DO <= x"00000000"; 
      when 3311 => DO <= x"00000000"; 
      when 3312 => DO <= x"00000000"; 
      when 3313 => DO <= x"00000000"; 
      when 3314 => DO <= x"00000000"; 
      when 3315 => DO <= x"00000000"; 
      when 3316 => DO <= x"00000000"; 
      when 3317 => DO <= x"00000000"; 
      when 3318 => DO <= x"00000000"; 
      when 3319 => DO <= x"00000000"; 
      when 3320 => DO <= x"00000000"; 
      when 3321 => DO <= x"00000000"; 
      when 3322 => DO <= x"00000000"; 
      when 3323 => DO <= x"00000000"; 
      when 3324 => DO <= x"00000000"; 
      when 3325 => DO <= x"00000000"; 
      when 3326 => DO <= x"00000000"; 
      when 3327 => DO <= x"00000000"; 
      when 3328 => DO <= x"00000000"; 
      when 3329 => DO <= x"00000000"; 
      when 3330 => DO <= x"00000000"; 
      when 3331 => DO <= x"00000000"; 
      when 3332 => DO <= x"00000000"; 
      when 3333 => DO <= x"00000000"; 
      when 3334 => DO <= x"00000000"; 
      when 3335 => DO <= x"00000000"; 
      when 3336 => DO <= x"00000000"; 
      when 3337 => DO <= x"00000000"; 
      when 3338 => DO <= x"00000000"; 
      when 3339 => DO <= x"00000000"; 
      when 3340 => DO <= x"00000000"; 
      when 3341 => DO <= x"00000000"; 
      when 3342 => DO <= x"00000000"; 
      when 3343 => DO <= x"00000000"; 
      when 3344 => DO <= x"00000000"; 
      when 3345 => DO <= x"00000000"; 
      when 3346 => DO <= x"00000000"; 
      when 3347 => DO <= x"00000000"; 
      when 3348 => DO <= x"00000000"; 
      when 3349 => DO <= x"00000000"; 
      when 3350 => DO <= x"00000000"; 
      when 3351 => DO <= x"00000000"; 
      when 3352 => DO <= x"00000000"; 
      when 3353 => DO <= x"00000000"; 
      when 3354 => DO <= x"00000000"; 
      when 3355 => DO <= x"00000000"; 
      when 3356 => DO <= x"00000000"; 
      when 3357 => DO <= x"00000000"; 
      when 3358 => DO <= x"00000000"; 
      when 3359 => DO <= x"00000000"; 
      when 3360 => DO <= x"00000000"; 
      when 3361 => DO <= x"00000000"; 
      when 3362 => DO <= x"00000000"; 
      when 3363 => DO <= x"00000000"; 
      when 3364 => DO <= x"00000000"; 
      when 3365 => DO <= x"00000000"; 
      when 3366 => DO <= x"00000000"; 
      when 3367 => DO <= x"00000000"; 
      when 3368 => DO <= x"00000000"; 
      when 3369 => DO <= x"00000000"; 
      when 3370 => DO <= x"00000000"; 
      when 3371 => DO <= x"00000000"; 
      when 3372 => DO <= x"00000000"; 
      when 3373 => DO <= x"00000000"; 
      when 3374 => DO <= x"00000000"; 
      when 3375 => DO <= x"00000000"; 
      when 3376 => DO <= x"00000000"; 
      when 3377 => DO <= x"00000000"; 
      when 3378 => DO <= x"00000000"; 
      when 3379 => DO <= x"00000000"; 
      when 3380 => DO <= x"00000000"; 
      when 3381 => DO <= x"00000000"; 
      when 3382 => DO <= x"00000000"; 
      when 3383 => DO <= x"00000000"; 
      when 3384 => DO <= x"00000000"; 
      when 3385 => DO <= x"00000000"; 
      when 3386 => DO <= x"00000000"; 
      when 3387 => DO <= x"00000000"; 
      when 3388 => DO <= x"00000000"; 
      when 3389 => DO <= x"00000000"; 
      when 3390 => DO <= x"00000000"; 
      when 3391 => DO <= x"00000000"; 
      when 3392 => DO <= x"00000000"; 
      when 3393 => DO <= x"00000000"; 
      when 3394 => DO <= x"00000000"; 
      when 3395 => DO <= x"00000000"; 
      when 3396 => DO <= x"00000000"; 
      when 3397 => DO <= x"00000000"; 
      when 3398 => DO <= x"00000000"; 
      when 3399 => DO <= x"00000000"; 
      when 3400 => DO <= x"00000000"; 
      when 3401 => DO <= x"00000000"; 
      when 3402 => DO <= x"00000000"; 
      when 3403 => DO <= x"00000000"; 
      when 3404 => DO <= x"00000000"; 
      when 3405 => DO <= x"00000000"; 
      when 3406 => DO <= x"00000000"; 
      when 3407 => DO <= x"00000000"; 
      when 3408 => DO <= x"00000000"; 
      when 3409 => DO <= x"00000000"; 
      when 3410 => DO <= x"00000000"; 
      when 3411 => DO <= x"00000000"; 
      when 3412 => DO <= x"00000000"; 
      when 3413 => DO <= x"00000000"; 
      when 3414 => DO <= x"00000000"; 
      when 3415 => DO <= x"00000000"; 
      when 3416 => DO <= x"00000000"; 
      when 3417 => DO <= x"00000000"; 
      when 3418 => DO <= x"00000000"; 
      when 3419 => DO <= x"00000000"; 
      when 3420 => DO <= x"00000000"; 
      when 3421 => DO <= x"00000000"; 
      when 3422 => DO <= x"00000000"; 
      when 3423 => DO <= x"00000000"; 
      when 3424 => DO <= x"00000000"; 
      when 3425 => DO <= x"00000000"; 
      when 3426 => DO <= x"00000000"; 
      when 3427 => DO <= x"00000000"; 
      when 3428 => DO <= x"00000000"; 
      when 3429 => DO <= x"00000000"; 
      when 3430 => DO <= x"00000000"; 
      when 3431 => DO <= x"00000000"; 
      when 3432 => DO <= x"00000000"; 
      when 3433 => DO <= x"00000000"; 
      when 3434 => DO <= x"00000000"; 
      when 3435 => DO <= x"00000000"; 
      when 3436 => DO <= x"00000000"; 
      when 3437 => DO <= x"00000000"; 
      when 3438 => DO <= x"00000000"; 
      when 3439 => DO <= x"00000000"; 
      when 3440 => DO <= x"00000000"; 
      when 3441 => DO <= x"00000000"; 
      when 3442 => DO <= x"00000000"; 
      when 3443 => DO <= x"00000000"; 
      when 3444 => DO <= x"00000000"; 
      when 3445 => DO <= x"00000000"; 
      when 3446 => DO <= x"00000000"; 
      when 3447 => DO <= x"00000000"; 
      when 3448 => DO <= x"00000000"; 
      when 3449 => DO <= x"00000000"; 
      when 3450 => DO <= x"00000000"; 
      when 3451 => DO <= x"00000000"; 
      when 3452 => DO <= x"00000000"; 
      when 3453 => DO <= x"00000000"; 
      when 3454 => DO <= x"00000000"; 
      when 3455 => DO <= x"00000000"; 
      when 3456 => DO <= x"00000000"; 
      when 3457 => DO <= x"00000000"; 
      when 3458 => DO <= x"00000000"; 
      when 3459 => DO <= x"00000000"; 
      when 3460 => DO <= x"00000000"; 
      when 3461 => DO <= x"00000000"; 
      when 3462 => DO <= x"00000000"; 
      when 3463 => DO <= x"00000000"; 
      when 3464 => DO <= x"00000000"; 
      when 3465 => DO <= x"00000000"; 
      when 3466 => DO <= x"00000000"; 
      when 3467 => DO <= x"00000000"; 
      when 3468 => DO <= x"00000000"; 
      when 3469 => DO <= x"00000000"; 
      when 3470 => DO <= x"00000000"; 
      when 3471 => DO <= x"00000000"; 
      when 3472 => DO <= x"00000000"; 
      when 3473 => DO <= x"00000000"; 
      when 3474 => DO <= x"00000000"; 
      when 3475 => DO <= x"00000000"; 
      when 3476 => DO <= x"00000000"; 
      when 3477 => DO <= x"00000000"; 
      when 3478 => DO <= x"00000000"; 
      when 3479 => DO <= x"00000000"; 
      when 3480 => DO <= x"00000000"; 
      when 3481 => DO <= x"00000000"; 
      when 3482 => DO <= x"00000000"; 
      when 3483 => DO <= x"00000000"; 
      when 3484 => DO <= x"00000000"; 
      when 3485 => DO <= x"00000000"; 
      when 3486 => DO <= x"00000000"; 
      when 3487 => DO <= x"00000000"; 
      when 3488 => DO <= x"00000000"; 
      when 3489 => DO <= x"00000000"; 
      when 3490 => DO <= x"00000000"; 
      when 3491 => DO <= x"00000000"; 
      when 3492 => DO <= x"00000000"; 
      when 3493 => DO <= x"00000000"; 
      when 3494 => DO <= x"00000000"; 
      when 3495 => DO <= x"00000000"; 
      when 3496 => DO <= x"00000000"; 
      when 3497 => DO <= x"00000000"; 
      when 3498 => DO <= x"00000000"; 
      when 3499 => DO <= x"00000000"; 
      when 3500 => DO <= x"00000000"; 
      when 3501 => DO <= x"00000000"; 
      when 3502 => DO <= x"00000000"; 
      when 3503 => DO <= x"00000000"; 
      when 3504 => DO <= x"00000000"; 
      when 3505 => DO <= x"00000000"; 
      when 3506 => DO <= x"00000000"; 
      when 3507 => DO <= x"00000000"; 
      when 3508 => DO <= x"00000000"; 
      when 3509 => DO <= x"00000000"; 
      when 3510 => DO <= x"00000000"; 
      when 3511 => DO <= x"00000000"; 
      when 3512 => DO <= x"00000000"; 
      when 3513 => DO <= x"00000000"; 
      when 3514 => DO <= x"00000000"; 
      when 3515 => DO <= x"00000000"; 
      when 3516 => DO <= x"00000000"; 
      when 3517 => DO <= x"00000000"; 
      when 3518 => DO <= x"00000000"; 
      when 3519 => DO <= x"00000000"; 
      when 3520 => DO <= x"00000000"; 
      when 3521 => DO <= x"00000000"; 
      when 3522 => DO <= x"00000000"; 
      when 3523 => DO <= x"00000000"; 
      when 3524 => DO <= x"00000000"; 
      when 3525 => DO <= x"00000000"; 
      when 3526 => DO <= x"00000000"; 
      when 3527 => DO <= x"00000000"; 
      when 3528 => DO <= x"00000000"; 
      when 3529 => DO <= x"00000000"; 
      when 3530 => DO <= x"00000000"; 
      when 3531 => DO <= x"00000000"; 
      when 3532 => DO <= x"00000000"; 
      when 3533 => DO <= x"00000000"; 
      when 3534 => DO <= x"00000000"; 
      when 3535 => DO <= x"00000000"; 
      when 3536 => DO <= x"00000000"; 
      when 3537 => DO <= x"00000000"; 
      when 3538 => DO <= x"00000000"; 
      when 3539 => DO <= x"00000000"; 
      when 3540 => DO <= x"00000000"; 
      when 3541 => DO <= x"00000000"; 
      when 3542 => DO <= x"00000000"; 
      when 3543 => DO <= x"00000000"; 
      when 3544 => DO <= x"00000000"; 
      when 3545 => DO <= x"00000000"; 
      when 3546 => DO <= x"00000000"; 
      when 3547 => DO <= x"00000000"; 
      when 3548 => DO <= x"00000000"; 
      when 3549 => DO <= x"00000000"; 
      when 3550 => DO <= x"00000000"; 
      when 3551 => DO <= x"00000000"; 
      when 3552 => DO <= x"00000000"; 
      when 3553 => DO <= x"00000000"; 
      when 3554 => DO <= x"00000000"; 
      when 3555 => DO <= x"00000000"; 
      when 3556 => DO <= x"00000000"; 
      when 3557 => DO <= x"00000000"; 
      when 3558 => DO <= x"00000000"; 
      when 3559 => DO <= x"00000000"; 
      when 3560 => DO <= x"00000000"; 
      when 3561 => DO <= x"00000000"; 
      when 3562 => DO <= x"00000000"; 
      when 3563 => DO <= x"00000000"; 
      when 3564 => DO <= x"00000000"; 
      when 3565 => DO <= x"00000000"; 
      when 3566 => DO <= x"00000000"; 
      when 3567 => DO <= x"00000000"; 
      when 3568 => DO <= x"00000000"; 
      when 3569 => DO <= x"00000000"; 
      when 3570 => DO <= x"00000000"; 
      when 3571 => DO <= x"00000000"; 
      when 3572 => DO <= x"00000000"; 
      when 3573 => DO <= x"00000000"; 
      when 3574 => DO <= x"00000000"; 
      when 3575 => DO <= x"00000000"; 
      when 3576 => DO <= x"00000000"; 
      when 3577 => DO <= x"00000000"; 
      when 3578 => DO <= x"00000000"; 
      when 3579 => DO <= x"00000000"; 
      when 3580 => DO <= x"00000000"; 
      when 3581 => DO <= x"00000000"; 
      when 3582 => DO <= x"00000000"; 
      when 3583 => DO <= x"00000000"; 
      when 3584 => DO <= x"00000000"; 
      when 3585 => DO <= x"00000000"; 
      when 3586 => DO <= x"00000000"; 
      when 3587 => DO <= x"00000000"; 
      when 3588 => DO <= x"00000000"; 
      when 3589 => DO <= x"00000000"; 
      when 3590 => DO <= x"00000000"; 
      when 3591 => DO <= x"00000000"; 
      when 3592 => DO <= x"00000000"; 
      when 3593 => DO <= x"00000000"; 
      when 3594 => DO <= x"00000000"; 
      when 3595 => DO <= x"00000000"; 
      when 3596 => DO <= x"00000000"; 
      when 3597 => DO <= x"00000000"; 
      when 3598 => DO <= x"00000000"; 
      when 3599 => DO <= x"00000000"; 
      when 3600 => DO <= x"00000000"; 
      when 3601 => DO <= x"00000000"; 
      when 3602 => DO <= x"00000000"; 
      when 3603 => DO <= x"00000000"; 
      when 3604 => DO <= x"00000000"; 
      when 3605 => DO <= x"00000000"; 
      when 3606 => DO <= x"00000000"; 
      when 3607 => DO <= x"00000000"; 
      when 3608 => DO <= x"00000000"; 
      when 3609 => DO <= x"00000000"; 
      when 3610 => DO <= x"00000000"; 
      when 3611 => DO <= x"00000000"; 
      when 3612 => DO <= x"00000000"; 
      when 3613 => DO <= x"00000000"; 
      when 3614 => DO <= x"00000000"; 
      when 3615 => DO <= x"00000000"; 
      when 3616 => DO <= x"00000000"; 
      when 3617 => DO <= x"00000000"; 
      when 3618 => DO <= x"00000000"; 
      when 3619 => DO <= x"00000000"; 
      when 3620 => DO <= x"00000000"; 
      when 3621 => DO <= x"00000000"; 
      when 3622 => DO <= x"00000000"; 
      when 3623 => DO <= x"00000000"; 
      when 3624 => DO <= x"00000000"; 
      when 3625 => DO <= x"00000000"; 
      when 3626 => DO <= x"00000000"; 
      when 3627 => DO <= x"00000000"; 
      when 3628 => DO <= x"00000000"; 
      when 3629 => DO <= x"00000000"; 
      when 3630 => DO <= x"00000000"; 
      when 3631 => DO <= x"00000000"; 
      when 3632 => DO <= x"00000000"; 
      when 3633 => DO <= x"00000000"; 
      when 3634 => DO <= x"00000000"; 
      when 3635 => DO <= x"00000000"; 
      when 3636 => DO <= x"00000000"; 
      when 3637 => DO <= x"00000000"; 
      when 3638 => DO <= x"00000000"; 
      when 3639 => DO <= x"00000000"; 
      when 3640 => DO <= x"00000000"; 
      when 3641 => DO <= x"00000000"; 
      when 3642 => DO <= x"00000000"; 
      when 3643 => DO <= x"00000000"; 
      when 3644 => DO <= x"00000000"; 
      when 3645 => DO <= x"00000000"; 
      when 3646 => DO <= x"00000000"; 
      when 3647 => DO <= x"00000000"; 
      when 3648 => DO <= x"00000000"; 
      when 3649 => DO <= x"00000000"; 
      when 3650 => DO <= x"00000000"; 
      when 3651 => DO <= x"00000000"; 
      when 3652 => DO <= x"00000000"; 
      when 3653 => DO <= x"00000000"; 
      when 3654 => DO <= x"00000000"; 
      when 3655 => DO <= x"00000000"; 
      when 3656 => DO <= x"00000000"; 
      when 3657 => DO <= x"00000000"; 
      when 3658 => DO <= x"00000000"; 
      when 3659 => DO <= x"00000000"; 
      when 3660 => DO <= x"00000000"; 
      when 3661 => DO <= x"00000000"; 
      when 3662 => DO <= x"00000000"; 
      when 3663 => DO <= x"00000000"; 
      when 3664 => DO <= x"00000000"; 
      when 3665 => DO <= x"00000000"; 
      when 3666 => DO <= x"00000000"; 
      when 3667 => DO <= x"00000000"; 
      when 3668 => DO <= x"00000000"; 
      when 3669 => DO <= x"00000000"; 
      when 3670 => DO <= x"00000000"; 
      when 3671 => DO <= x"00000000"; 
      when 3672 => DO <= x"00000000"; 
      when 3673 => DO <= x"00000000"; 
      when 3674 => DO <= x"00000000"; 
      when 3675 => DO <= x"00000000"; 
      when 3676 => DO <= x"00000000"; 
      when 3677 => DO <= x"00000000"; 
      when 3678 => DO <= x"00000000"; 
      when 3679 => DO <= x"00000000"; 
      when 3680 => DO <= x"00000000"; 
      when 3681 => DO <= x"00000000"; 
      when 3682 => DO <= x"00000000"; 
      when 3683 => DO <= x"00000000"; 
      when 3684 => DO <= x"00000000"; 
      when 3685 => DO <= x"00000000"; 
      when 3686 => DO <= x"00000000"; 
      when 3687 => DO <= x"00000000"; 
      when 3688 => DO <= x"00000000"; 
      when 3689 => DO <= x"00000000"; 
      when 3690 => DO <= x"00000000"; 
      when 3691 => DO <= x"00000000"; 
      when 3692 => DO <= x"00000000"; 
      when 3693 => DO <= x"00000000"; 
      when 3694 => DO <= x"00000000"; 
      when 3695 => DO <= x"00000000"; 
      when 3696 => DO <= x"00000000"; 
      when 3697 => DO <= x"00000000"; 
      when 3698 => DO <= x"00000000"; 
      when 3699 => DO <= x"00000000"; 
      when 3700 => DO <= x"00000000"; 
      when 3701 => DO <= x"00000000"; 
      when 3702 => DO <= x"00000000"; 
      when 3703 => DO <= x"00000000"; 
      when 3704 => DO <= x"00000000"; 
      when 3705 => DO <= x"00000000"; 
      when 3706 => DO <= x"00000000"; 
      when 3707 => DO <= x"00000000"; 
      when 3708 => DO <= x"00000000"; 
      when 3709 => DO <= x"00000000"; 
      when 3710 => DO <= x"00000000"; 
      when 3711 => DO <= x"00000000"; 
      when 3712 => DO <= x"00000000"; 
      when 3713 => DO <= x"00000000"; 
      when 3714 => DO <= x"00000000"; 
      when 3715 => DO <= x"00000000"; 
      when 3716 => DO <= x"00000000"; 
      when 3717 => DO <= x"00000000"; 
      when 3718 => DO <= x"00000000"; 
      when 3719 => DO <= x"00000000"; 
      when 3720 => DO <= x"00000000"; 
      when 3721 => DO <= x"00000000"; 
      when 3722 => DO <= x"00000000"; 
      when 3723 => DO <= x"00000000"; 
      when 3724 => DO <= x"00000000"; 
      when 3725 => DO <= x"00000000"; 
      when 3726 => DO <= x"00000000"; 
      when 3727 => DO <= x"00000000"; 
      when 3728 => DO <= x"00000000"; 
      when 3729 => DO <= x"00000000"; 
      when 3730 => DO <= x"00000000"; 
      when 3731 => DO <= x"00000000"; 
      when 3732 => DO <= x"00000000"; 
      when 3733 => DO <= x"00000000"; 
      when 3734 => DO <= x"00000000"; 
      when 3735 => DO <= x"00000000"; 
      when 3736 => DO <= x"00000000"; 
      when 3737 => DO <= x"00000000"; 
      when 3738 => DO <= x"00000000"; 
      when 3739 => DO <= x"00000000"; 
      when 3740 => DO <= x"00000000"; 
      when 3741 => DO <= x"00000000"; 
      when 3742 => DO <= x"00000000"; 
      when 3743 => DO <= x"00000000"; 
      when 3744 => DO <= x"00000000"; 
      when 3745 => DO <= x"00000000"; 
      when 3746 => DO <= x"00000000"; 
      when 3747 => DO <= x"00000000"; 
      when 3748 => DO <= x"00000000"; 
      when 3749 => DO <= x"00000000"; 
      when 3750 => DO <= x"00000000"; 
      when 3751 => DO <= x"00000000"; 
      when 3752 => DO <= x"00000000"; 
      when 3753 => DO <= x"00000000"; 
      when 3754 => DO <= x"00000000"; 
      when 3755 => DO <= x"00000000"; 
      when 3756 => DO <= x"00000000"; 
      when 3757 => DO <= x"00000000"; 
      when 3758 => DO <= x"00000000"; 
      when 3759 => DO <= x"00000000"; 
      when 3760 => DO <= x"00000000"; 
      when 3761 => DO <= x"00000000"; 
      when 3762 => DO <= x"00000000"; 
      when 3763 => DO <= x"00000000"; 
      when 3764 => DO <= x"00000000"; 
      when 3765 => DO <= x"00000000"; 
      when 3766 => DO <= x"00000000"; 
      when 3767 => DO <= x"00000000"; 
      when 3768 => DO <= x"00000000"; 
      when 3769 => DO <= x"00000000"; 
      when 3770 => DO <= x"00000000"; 
      when 3771 => DO <= x"00000000"; 
      when 3772 => DO <= x"00000000"; 
      when 3773 => DO <= x"00000000"; 
      when 3774 => DO <= x"00000000"; 
      when 3775 => DO <= x"00000000"; 
      when 3776 => DO <= x"00000000"; 
      when 3777 => DO <= x"00000000"; 
      when 3778 => DO <= x"00000000"; 
      when 3779 => DO <= x"00000000"; 
      when 3780 => DO <= x"00000000"; 
      when 3781 => DO <= x"00000000"; 
      when 3782 => DO <= x"00000000"; 
      when 3783 => DO <= x"00000000"; 
      when 3784 => DO <= x"00000000"; 
      when 3785 => DO <= x"00000000"; 
      when 3786 => DO <= x"00000000"; 
      when 3787 => DO <= x"00000000"; 
      when 3788 => DO <= x"00000000"; 
      when 3789 => DO <= x"00000000"; 
      when 3790 => DO <= x"00000000"; 
      when 3791 => DO <= x"00000000"; 
      when 3792 => DO <= x"00000000"; 
      when 3793 => DO <= x"00000000"; 
      when 3794 => DO <= x"00000000"; 
      when 3795 => DO <= x"00000000"; 
      when 3796 => DO <= x"00000000"; 
      when 3797 => DO <= x"00000000"; 
      when 3798 => DO <= x"00000000"; 
      when 3799 => DO <= x"00000000"; 
      when 3800 => DO <= x"00000000"; 
      when 3801 => DO <= x"00000000"; 
      when 3802 => DO <= x"00000000"; 
      when 3803 => DO <= x"00000000"; 
      when 3804 => DO <= x"00000000"; 
      when 3805 => DO <= x"00000000"; 
      when 3806 => DO <= x"00000000"; 
      when 3807 => DO <= x"00000000"; 
      when 3808 => DO <= x"00000000"; 
      when 3809 => DO <= x"00000000"; 
      when 3810 => DO <= x"00000000"; 
      when 3811 => DO <= x"00000000"; 
      when 3812 => DO <= x"00000000"; 
      when 3813 => DO <= x"00000000"; 
      when 3814 => DO <= x"00000000"; 
      when 3815 => DO <= x"00000000"; 
      when 3816 => DO <= x"00000000"; 
      when 3817 => DO <= x"00000000"; 
      when 3818 => DO <= x"00000000"; 
      when 3819 => DO <= x"00000000"; 
      when 3820 => DO <= x"00000000"; 
      when 3821 => DO <= x"00000000"; 
      when 3822 => DO <= x"00000000"; 
      when 3823 => DO <= x"00000000"; 
      when 3824 => DO <= x"00000000"; 
      when 3825 => DO <= x"00000000"; 
      when 3826 => DO <= x"00000000"; 
      when 3827 => DO <= x"00000000"; 
      when 3828 => DO <= x"00000000"; 
      when 3829 => DO <= x"00000000"; 
      when 3830 => DO <= x"00000000"; 
      when 3831 => DO <= x"00000000"; 
      when 3832 => DO <= x"00000000"; 
      when 3833 => DO <= x"00000000"; 
      when 3834 => DO <= x"00000000"; 
      when 3835 => DO <= x"00000000"; 
      when 3836 => DO <= x"00000000"; 
      when 3837 => DO <= x"00000000"; 
      when 3838 => DO <= x"00000000"; 
      when 3839 => DO <= x"00000000"; 
      when 3840 => DO <= x"00000000"; 
      when 3841 => DO <= x"00000000"; 
      when 3842 => DO <= x"00000000"; 
      when 3843 => DO <= x"00000000"; 
      when 3844 => DO <= x"00000000"; 
      when 3845 => DO <= x"00000000"; 
      when 3846 => DO <= x"00000000"; 
      when 3847 => DO <= x"00000000"; 
      when 3848 => DO <= x"00000000"; 
      when 3849 => DO <= x"00000000"; 
      when 3850 => DO <= x"00000000"; 
      when 3851 => DO <= x"00000000"; 
      when 3852 => DO <= x"00000000"; 
      when 3853 => DO <= x"00000000"; 
      when 3854 => DO <= x"00000000"; 
      when 3855 => DO <= x"00000000"; 
      when 3856 => DO <= x"00000000"; 
      when 3857 => DO <= x"00000000"; 
      when 3858 => DO <= x"00000000"; 
      when 3859 => DO <= x"00000000"; 
      when 3860 => DO <= x"00000000"; 
      when 3861 => DO <= x"00000000"; 
      when 3862 => DO <= x"00000000"; 
      when 3863 => DO <= x"00000000"; 
      when 3864 => DO <= x"00000000"; 
      when 3865 => DO <= x"00000000"; 
      when 3866 => DO <= x"00000000"; 
      when 3867 => DO <= x"00000000"; 
      when 3868 => DO <= x"00000000"; 
      when 3869 => DO <= x"00000000"; 
      when 3870 => DO <= x"00000000"; 
      when 3871 => DO <= x"00000000"; 
      when 3872 => DO <= x"00000000"; 
      when 3873 => DO <= x"00000000"; 
      when 3874 => DO <= x"00000000"; 
      when 3875 => DO <= x"00000000"; 
      when 3876 => DO <= x"00000000"; 
      when 3877 => DO <= x"00000000"; 
      when 3878 => DO <= x"00000000"; 
      when 3879 => DO <= x"00000000"; 
      when 3880 => DO <= x"00000000"; 
      when 3881 => DO <= x"00000000"; 
      when 3882 => DO <= x"00000000"; 
      when 3883 => DO <= x"00000000"; 
      when 3884 => DO <= x"00000000"; 
      when 3885 => DO <= x"00000000"; 
      when 3886 => DO <= x"00000000"; 
      when 3887 => DO <= x"00000000"; 
      when 3888 => DO <= x"00000000"; 
      when 3889 => DO <= x"00000000"; 
      when 3890 => DO <= x"00000000"; 
      when 3891 => DO <= x"00000000"; 
      when 3892 => DO <= x"00000000"; 
      when 3893 => DO <= x"00000000"; 
      when 3894 => DO <= x"00000000"; 
      when 3895 => DO <= x"00000000"; 
      when 3896 => DO <= x"00000000"; 
      when 3897 => DO <= x"00000000"; 
      when 3898 => DO <= x"00000000"; 
      when 3899 => DO <= x"00000000"; 
      when 3900 => DO <= x"00000000"; 
      when 3901 => DO <= x"00000000"; 
      when 3902 => DO <= x"00000000"; 
      when 3903 => DO <= x"00000000"; 
      when 3904 => DO <= x"00000000"; 
      when 3905 => DO <= x"00000000"; 
      when 3906 => DO <= x"00000000"; 
      when 3907 => DO <= x"00000000"; 
      when 3908 => DO <= x"00000000"; 
      when 3909 => DO <= x"00000000"; 
      when 3910 => DO <= x"00000000"; 
      when 3911 => DO <= x"00000000"; 
      when 3912 => DO <= x"00000000"; 
      when 3913 => DO <= x"00000000"; 
      when 3914 => DO <= x"00000000"; 
      when 3915 => DO <= x"00000000"; 
      when 3916 => DO <= x"00000000"; 
      when 3917 => DO <= x"00000000"; 
      when 3918 => DO <= x"00000000"; 
      when 3919 => DO <= x"00000000"; 
      when 3920 => DO <= x"00000000"; 
      when 3921 => DO <= x"00000000"; 
      when 3922 => DO <= x"00000000"; 
      when 3923 => DO <= x"00000000"; 
      when 3924 => DO <= x"00000000"; 
      when 3925 => DO <= x"00000000"; 
      when 3926 => DO <= x"00000000"; 
      when 3927 => DO <= x"00000000"; 
      when 3928 => DO <= x"00000000"; 
      when 3929 => DO <= x"00000000"; 
      when 3930 => DO <= x"00000000"; 
      when 3931 => DO <= x"00000000"; 
      when 3932 => DO <= x"00000000"; 
      when 3933 => DO <= x"00000000"; 
      when 3934 => DO <= x"00000000"; 
      when 3935 => DO <= x"00000000"; 
      when 3936 => DO <= x"00000000"; 
      when 3937 => DO <= x"00000000"; 
      when 3938 => DO <= x"00000000"; 
      when 3939 => DO <= x"00000000"; 
      when 3940 => DO <= x"00000000"; 
      when 3941 => DO <= x"00000000"; 
      when 3942 => DO <= x"00000000"; 
      when 3943 => DO <= x"00000000"; 
      when 3944 => DO <= x"00000000"; 
      when 3945 => DO <= x"00000000"; 
      when 3946 => DO <= x"00000000"; 
      when 3947 => DO <= x"00000000"; 
      when 3948 => DO <= x"00000000"; 
      when 3949 => DO <= x"00000000"; 
      when 3950 => DO <= x"00000000"; 
      when 3951 => DO <= x"00000000"; 
      when 3952 => DO <= x"00000000"; 
      when 3953 => DO <= x"00000000"; 
      when 3954 => DO <= x"00000000"; 
      when 3955 => DO <= x"00000000"; 
      when 3956 => DO <= x"00000000"; 
      when 3957 => DO <= x"00000000"; 
      when 3958 => DO <= x"00000000"; 
      when 3959 => DO <= x"00000000"; 
      when 3960 => DO <= x"00000000"; 
      when 3961 => DO <= x"00000000"; 
      when 3962 => DO <= x"00000000"; 
      when 3963 => DO <= x"00000000"; 
      when 3964 => DO <= x"00000000"; 
      when 3965 => DO <= x"00000000"; 
      when 3966 => DO <= x"00000000"; 
      when 3967 => DO <= x"00000000"; 
      when 3968 => DO <= x"00000000"; 
      when 3969 => DO <= x"00000000"; 
      when 3970 => DO <= x"00000000"; 
      when 3971 => DO <= x"00000000"; 
      when 3972 => DO <= x"00000000"; 
      when 3973 => DO <= x"00000000"; 
      when 3974 => DO <= x"00000000"; 
      when 3975 => DO <= x"00000000"; 
      when 3976 => DO <= x"00000000"; 
      when 3977 => DO <= x"00000000"; 
      when 3978 => DO <= x"00000000"; 
      when 3979 => DO <= x"00000000"; 
      when 3980 => DO <= x"00000000"; 
      when 3981 => DO <= x"00000000"; 
      when 3982 => DO <= x"00000000"; 
      when 3983 => DO <= x"00000000"; 
      when 3984 => DO <= x"00000000"; 
      when 3985 => DO <= x"00000000"; 
      when 3986 => DO <= x"00000000"; 
      when 3987 => DO <= x"00000000"; 
      when 3988 => DO <= x"00000000"; 
      when 3989 => DO <= x"00000000"; 
      when 3990 => DO <= x"00000000"; 
      when 3991 => DO <= x"00000000"; 
      when 3992 => DO <= x"00000000"; 
      when 3993 => DO <= x"00000000"; 
      when 3994 => DO <= x"00000000"; 
      when 3995 => DO <= x"00000000"; 
      when 3996 => DO <= x"00000000"; 
      when 3997 => DO <= x"00000000"; 
      when 3998 => DO <= x"00000000"; 
      when 3999 => DO <= x"00000000"; 
      when 4000 => DO <= x"00000000"; 
      when 4001 => DO <= x"00000000"; 
      when 4002 => DO <= x"00000000"; 
      when 4003 => DO <= x"00000000"; 
      when 4004 => DO <= x"00000000"; 
      when 4005 => DO <= x"00000000"; 
      when 4006 => DO <= x"00000000"; 
      when 4007 => DO <= x"00000000"; 
      when 4008 => DO <= x"00000000"; 
      when 4009 => DO <= x"00000000"; 
      when 4010 => DO <= x"00000000"; 
      when 4011 => DO <= x"00000000"; 
      when 4012 => DO <= x"00000000"; 
      when 4013 => DO <= x"00000000"; 
      when 4014 => DO <= x"00000000"; 
      when 4015 => DO <= x"00000000"; 
      when 4016 => DO <= x"00000000"; 
      when 4017 => DO <= x"00000000"; 
      when 4018 => DO <= x"00000000"; 
      when 4019 => DO <= x"00000000"; 
      when 4020 => DO <= x"00000000"; 
      when 4021 => DO <= x"00000000"; 
      when 4022 => DO <= x"00000000"; 
      when 4023 => DO <= x"00000000"; 
      when 4024 => DO <= x"00000000"; 
      when 4025 => DO <= x"00000000"; 
      when 4026 => DO <= x"00000000"; 
      when 4027 => DO <= x"00000000"; 
      when 4028 => DO <= x"00000000"; 
      when 4029 => DO <= x"00000000"; 
      when 4030 => DO <= x"00000000"; 
      when 4031 => DO <= x"00000000"; 
      when 4032 => DO <= x"00000000"; 
      when 4033 => DO <= x"00000000"; 
      when 4034 => DO <= x"00000000"; 
      when 4035 => DO <= x"00000000"; 
      when 4036 => DO <= x"00000000"; 
      when 4037 => DO <= x"00000000"; 
      when 4038 => DO <= x"00000000"; 
      when 4039 => DO <= x"00000000"; 
      when 4040 => DO <= x"00000000"; 
      when 4041 => DO <= x"00000000"; 
      when 4042 => DO <= x"00000000"; 
      when 4043 => DO <= x"00000000"; 
      when 4044 => DO <= x"00000000"; 
      when 4045 => DO <= x"00000000"; 
      when 4046 => DO <= x"00000000"; 
      when 4047 => DO <= x"00000000"; 
      when 4048 => DO <= x"00000000"; 
      when 4049 => DO <= x"00000000"; 
      when 4050 => DO <= x"00000000"; 
      when 4051 => DO <= x"00000000"; 
      when 4052 => DO <= x"00000000"; 
      when 4053 => DO <= x"00000000"; 
      when 4054 => DO <= x"00000000"; 
      when 4055 => DO <= x"00000000"; 
      when 4056 => DO <= x"00000000"; 
      when 4057 => DO <= x"00000000"; 
      when 4058 => DO <= x"00000000"; 
      when 4059 => DO <= x"00000000"; 
      when 4060 => DO <= x"00000000"; 
      when 4061 => DO <= x"00000000"; 
      when 4062 => DO <= x"00000000"; 
      when 4063 => DO <= x"00000000"; 
      when 4064 => DO <= x"00000000"; 
      when 4065 => DO <= x"00000000"; 
      when 4066 => DO <= x"00000000"; 
      when 4067 => DO <= x"00000000"; 
      when 4068 => DO <= x"00000000"; 
      when 4069 => DO <= x"00000000"; 
      when 4070 => DO <= x"00000000"; 
      when 4071 => DO <= x"00000000"; 
      when 4072 => DO <= x"00000000"; 
      when 4073 => DO <= x"00000000"; 
      when 4074 => DO <= x"00000000"; 
      when 4075 => DO <= x"00000000"; 
      when 4076 => DO <= x"00000000"; 
      when 4077 => DO <= x"00000000"; 
      when 4078 => DO <= x"00000000"; 
      when 4079 => DO <= x"00000000"; 
      when 4080 => DO <= x"00000000"; 
      when 4081 => DO <= x"00000000"; 
      when 4082 => DO <= x"00000000"; 
      when 4083 => DO <= x"00000000"; 
      when 4084 => DO <= x"00000000"; 
      when 4085 => DO <= x"00000000"; 
      when 4086 => DO <= x"00000000"; 
      when 4087 => DO <= x"00000000"; 
      when 4088 => DO <= x"00000000"; 
      when 4089 => DO <= x"00000000"; 
      when 4090 => DO <= x"00000000"; 
      when 4091 => DO <= x"00000000"; 
      when 4092 => DO <= x"00000000"; 
      when 4093 => DO <= x"00000000"; 
      when 4094 => DO <= x"00000000"; 
      when 4095 => DO <= x"00000000"; 
      when 4096 => DO <= x"00000000"; 
      when 4097 => DO <= x"00000000"; 
      when 4098 => DO <= x"00000000"; 
      when 4099 => DO <= x"00000000"; 
      when 4100 => DO <= x"00000000"; 
      when 4101 => DO <= x"00000000"; 
      when 4102 => DO <= x"00000000"; 
      when 4103 => DO <= x"00000000"; 
      when 4104 => DO <= x"00000000"; 
      when 4105 => DO <= x"00000000"; 
      when 4106 => DO <= x"00000000"; 
      when 4107 => DO <= x"00000000"; 
      when 4108 => DO <= x"00000000"; 
      when 4109 => DO <= x"00000000"; 
      when 4110 => DO <= x"00000000"; 
      when 4111 => DO <= x"00000000"; 
      when 4112 => DO <= x"00000000"; 
      when 4113 => DO <= x"00000000"; 
      when 4114 => DO <= x"00000000"; 
      when 4115 => DO <= x"00000000"; 
      when 4116 => DO <= x"00000000"; 
      when 4117 => DO <= x"00000000"; 
      when 4118 => DO <= x"00000000"; 
      when 4119 => DO <= x"00000000"; 
      when 4120 => DO <= x"00000000"; 
      when 4121 => DO <= x"00000000"; 
      when 4122 => DO <= x"00000000"; 
      when 4123 => DO <= x"00000000"; 
      when 4124 => DO <= x"00000000"; 
      when 4125 => DO <= x"00000000"; 
      when 4126 => DO <= x"00000000"; 
      when 4127 => DO <= x"00000000"; 
      when 4128 => DO <= x"00000000"; 
      when 4129 => DO <= x"00000000"; 
      when 4130 => DO <= x"00000000"; 
      when 4131 => DO <= x"00000000"; 
      when 4132 => DO <= x"00000000"; 
      when 4133 => DO <= x"00000000"; 
      when 4134 => DO <= x"00000000"; 
      when 4135 => DO <= x"00000000"; 
      when 4136 => DO <= x"00000000"; 
      when 4137 => DO <= x"00000000"; 
      when 4138 => DO <= x"00000000"; 
      when 4139 => DO <= x"00000000"; 
      when 4140 => DO <= x"00000000"; 
      when 4141 => DO <= x"00000000"; 
      when 4142 => DO <= x"00000000"; 
      when 4143 => DO <= x"00000000"; 
      when 4144 => DO <= x"00000000"; 
      when 4145 => DO <= x"00000000"; 
      when 4146 => DO <= x"00000000"; 
      when 4147 => DO <= x"00000000"; 
      when 4148 => DO <= x"00000000"; 
      when 4149 => DO <= x"00000000"; 
      when 4150 => DO <= x"00000000"; 
      when 4151 => DO <= x"00000000"; 
      when 4152 => DO <= x"00000000"; 
      when 4153 => DO <= x"00000000"; 
      when 4154 => DO <= x"00000000"; 
      when 4155 => DO <= x"00000000"; 
      when 4156 => DO <= x"00000000"; 
      when 4157 => DO <= x"00000000"; 
      when 4158 => DO <= x"00000000"; 
      when 4159 => DO <= x"00000000"; 
      when 4160 => DO <= x"00000000"; 
      when 4161 => DO <= x"00000000"; 
      when 4162 => DO <= x"00000000"; 
      when 4163 => DO <= x"00000000"; 
      when 4164 => DO <= x"00000000"; 
      when 4165 => DO <= x"00000000"; 
      when 4166 => DO <= x"00000000"; 
      when 4167 => DO <= x"00000000"; 
      when 4168 => DO <= x"00000000"; 
      when 4169 => DO <= x"00000000"; 
      when 4170 => DO <= x"00000000"; 
      when 4171 => DO <= x"00000000"; 
      when 4172 => DO <= x"00000000"; 
      when 4173 => DO <= x"00000000"; 
      when 4174 => DO <= x"00000000"; 
      when 4175 => DO <= x"00000000"; 
      when 4176 => DO <= x"00000000"; 
      when 4177 => DO <= x"00000000"; 
      when 4178 => DO <= x"00000000"; 
      when 4179 => DO <= x"00000000"; 
      when 4180 => DO <= x"00000000"; 
      when 4181 => DO <= x"00000000"; 
      when 4182 => DO <= x"00000000"; 
      when 4183 => DO <= x"00000000"; 
      when 4184 => DO <= x"00000000"; 
      when 4185 => DO <= x"00000000"; 
      when 4186 => DO <= x"00000000"; 
      when 4187 => DO <= x"00000000"; 
      when 4188 => DO <= x"00000000"; 
      when 4189 => DO <= x"00000000"; 
      when 4190 => DO <= x"00000000"; 
      when 4191 => DO <= x"00000000"; 
      when 4192 => DO <= x"00000000"; 
      when 4193 => DO <= x"00000000"; 
      when 4194 => DO <= x"00000000"; 
      when 4195 => DO <= x"00000000"; 
      when 4196 => DO <= x"00000000"; 
      when 4197 => DO <= x"00000000"; 
      when 4198 => DO <= x"00000000"; 
      when 4199 => DO <= x"00000000"; 
      when 4200 => DO <= x"00000000"; 
      when 4201 => DO <= x"00000000"; 
      when 4202 => DO <= x"00000000"; 
      when 4203 => DO <= x"00000000"; 
      when 4204 => DO <= x"00000000"; 
      when 4205 => DO <= x"00000000"; 
      when 4206 => DO <= x"00000000"; 
      when 4207 => DO <= x"00000000"; 
      when 4208 => DO <= x"00000000"; 
      when 4209 => DO <= x"00000000"; 
      when 4210 => DO <= x"00000000"; 
      when 4211 => DO <= x"00000000"; 
      when 4212 => DO <= x"00000000"; 
      when 4213 => DO <= x"00000000"; 
      when 4214 => DO <= x"00000000"; 
      when 4215 => DO <= x"00000000"; 
      when 4216 => DO <= x"00000000"; 
      when 4217 => DO <= x"00000000"; 
      when 4218 => DO <= x"00000000"; 
      when 4219 => DO <= x"00000000"; 
      when 4220 => DO <= x"00000000"; 
      when 4221 => DO <= x"00000000"; 
      when 4222 => DO <= x"00000000"; 
      when 4223 => DO <= x"00000000"; 
      when 4224 => DO <= x"00000000"; 
      when 4225 => DO <= x"00000000"; 
      when 4226 => DO <= x"00000000"; 
      when 4227 => DO <= x"00000000"; 
      when 4228 => DO <= x"00000000"; 
      when 4229 => DO <= x"00000000"; 
      when 4230 => DO <= x"00000000"; 
      when 4231 => DO <= x"00000000"; 
      when 4232 => DO <= x"00000000"; 
      when 4233 => DO <= x"00000000"; 
      when 4234 => DO <= x"00000000"; 
      when 4235 => DO <= x"00000000"; 
      when 4236 => DO <= x"00000000"; 
      when 4237 => DO <= x"00000000"; 
      when 4238 => DO <= x"00000000"; 
      when 4239 => DO <= x"00000000"; 
      when 4240 => DO <= x"00000000"; 
      when 4241 => DO <= x"00000000"; 
      when 4242 => DO <= x"00000000"; 
      when 4243 => DO <= x"00000000"; 
      when 4244 => DO <= x"00000000"; 
      when 4245 => DO <= x"00000000"; 
      when 4246 => DO <= x"00000000"; 
      when 4247 => DO <= x"00000000"; 
      when 4248 => DO <= x"00000000"; 
      when 4249 => DO <= x"00000000"; 
      when 4250 => DO <= x"00000000"; 
      when 4251 => DO <= x"00000000"; 
      when 4252 => DO <= x"00000000"; 
      when 4253 => DO <= x"00000000"; 
      when 4254 => DO <= x"00000000"; 
      when 4255 => DO <= x"00000000"; 
      when 4256 => DO <= x"00000000"; 
      when 4257 => DO <= x"00000000"; 
      when 4258 => DO <= x"00000000"; 
      when 4259 => DO <= x"00000000"; 
      when 4260 => DO <= x"00000000"; 
      when 4261 => DO <= x"00000000"; 
      when 4262 => DO <= x"00000000"; 
      when 4263 => DO <= x"00000000"; 
      when 4264 => DO <= x"00000000"; 
      when 4265 => DO <= x"00000000"; 
      when 4266 => DO <= x"00000000"; 
      when 4267 => DO <= x"00000000"; 
      when 4268 => DO <= x"00000000"; 
      when 4269 => DO <= x"00000000"; 
      when 4270 => DO <= x"00000000"; 
      when 4271 => DO <= x"00000000"; 
      when 4272 => DO <= x"00000000"; 
      when 4273 => DO <= x"00000000"; 
      when 4274 => DO <= x"00000000"; 
      when 4275 => DO <= x"00000000"; 
      when 4276 => DO <= x"00000000"; 
      when 4277 => DO <= x"00000000"; 
      when 4278 => DO <= x"00000000"; 
      when 4279 => DO <= x"00000000"; 
      when 4280 => DO <= x"00000000"; 
      when 4281 => DO <= x"00000000"; 
      when 4282 => DO <= x"00000000"; 
      when 4283 => DO <= x"00000000"; 
      when 4284 => DO <= x"00000000"; 
      when 4285 => DO <= x"00000000"; 
      when 4286 => DO <= x"00000000"; 
      when 4287 => DO <= x"00000000"; 
      when 4288 => DO <= x"00000000"; 
      when 4289 => DO <= x"00000000"; 
      when 4290 => DO <= x"00000000"; 
      when 4291 => DO <= x"00000000"; 
      when 4292 => DO <= x"00000000"; 
      when 4293 => DO <= x"00000000"; 
      when 4294 => DO <= x"00000000"; 
      when 4295 => DO <= x"00000000"; 
      when 4296 => DO <= x"00000000"; 
      when 4297 => DO <= x"00000000"; 
      when 4298 => DO <= x"00000000"; 
      when 4299 => DO <= x"00000000"; 
      when 4300 => DO <= x"00000000"; 
      when 4301 => DO <= x"00000000"; 
      when 4302 => DO <= x"00000000"; 
      when 4303 => DO <= x"00000000"; 
      when 4304 => DO <= x"00000000"; 
      when 4305 => DO <= x"00000000"; 
      when 4306 => DO <= x"00000000"; 
      when 4307 => DO <= x"00000000"; 
      when 4308 => DO <= x"00000000"; 
      when 4309 => DO <= x"00000000"; 
      when 4310 => DO <= x"00000000"; 
      when 4311 => DO <= x"00000000"; 
      when 4312 => DO <= x"00000000"; 
      when 4313 => DO <= x"00000000"; 
      when 4314 => DO <= x"00000000"; 
      when 4315 => DO <= x"00000000"; 
      when 4316 => DO <= x"00000000"; 
      when 4317 => DO <= x"00000000"; 
      when 4318 => DO <= x"00000000"; 
      when 4319 => DO <= x"00000000"; 
      when 4320 => DO <= x"00000000"; 
      when 4321 => DO <= x"00000000"; 
      when 4322 => DO <= x"00000000"; 
      when 4323 => DO <= x"00000000"; 
      when 4324 => DO <= x"00000000"; 
      when 4325 => DO <= x"00000000"; 
      when 4326 => DO <= x"00000000"; 
      when 4327 => DO <= x"00000000"; 
      when 4328 => DO <= x"00000000"; 
      when 4329 => DO <= x"00000000"; 
      when 4330 => DO <= x"00000000"; 
      when 4331 => DO <= x"00000000"; 
      when 4332 => DO <= x"00000000"; 
      when 4333 => DO <= x"00000000"; 
      when 4334 => DO <= x"00000000"; 
      when 4335 => DO <= x"00000000"; 
      when 4336 => DO <= x"00000000"; 
      when 4337 => DO <= x"00000000"; 
      when 4338 => DO <= x"00000000"; 
      when 4339 => DO <= x"00000000"; 
      when 4340 => DO <= x"00000000"; 
      when 4341 => DO <= x"00000000"; 
      when 4342 => DO <= x"00000000"; 
      when 4343 => DO <= x"00000000"; 
      when 4344 => DO <= x"00000000"; 
      when 4345 => DO <= x"00000000"; 
      when 4346 => DO <= x"00000000"; 
      when 4347 => DO <= x"00000000"; 
      when 4348 => DO <= x"00000000"; 
      when 4349 => DO <= x"00000000"; 
      when 4350 => DO <= x"00000000"; 
      when 4351 => DO <= x"00000000"; 
      when 4352 => DO <= x"00000000"; 
      when 4353 => DO <= x"00000000"; 
      when 4354 => DO <= x"00000000"; 
      when 4355 => DO <= x"00000000"; 
      when 4356 => DO <= x"00000000"; 
      when 4357 => DO <= x"00000000"; 
      when 4358 => DO <= x"00000000"; 
      when 4359 => DO <= x"00000000"; 
      when 4360 => DO <= x"00000000"; 
      when 4361 => DO <= x"00000000"; 
      when 4362 => DO <= x"00000000"; 
      when 4363 => DO <= x"00000000"; 
      when 4364 => DO <= x"00000000"; 
      when 4365 => DO <= x"00000000"; 
      when 4366 => DO <= x"00000000"; 
      when 4367 => DO <= x"00000000"; 
      when 4368 => DO <= x"00000000"; 
      when 4369 => DO <= x"00000000"; 
      when 4370 => DO <= x"00000000"; 
      when 4371 => DO <= x"00000000"; 
      when 4372 => DO <= x"00000000"; 
      when 4373 => DO <= x"00000000"; 
      when 4374 => DO <= x"00000000"; 
      when 4375 => DO <= x"00000000"; 
      when 4376 => DO <= x"00000000"; 
      when 4377 => DO <= x"00000000"; 
      when 4378 => DO <= x"00000000"; 
      when 4379 => DO <= x"00000000"; 
      when 4380 => DO <= x"00000000"; 
      when 4381 => DO <= x"00000000"; 
      when 4382 => DO <= x"00000000"; 
      when 4383 => DO <= x"00000000"; 
      when 4384 => DO <= x"00000000"; 
      when 4385 => DO <= x"00000000"; 
      when 4386 => DO <= x"00000000"; 
      when 4387 => DO <= x"00000000"; 
      when 4388 => DO <= x"00000000"; 
      when 4389 => DO <= x"00000000"; 
      when 4390 => DO <= x"00000000"; 
      when 4391 => DO <= x"00000000"; 
      when 4392 => DO <= x"00000000"; 
      when 4393 => DO <= x"00000000"; 
      when 4394 => DO <= x"00000000"; 
      when 4395 => DO <= x"00000000"; 
      when 4396 => DO <= x"00000000"; 
      when 4397 => DO <= x"00000000"; 
      when 4398 => DO <= x"00000000"; 
      when 4399 => DO <= x"00000000"; 
      when 4400 => DO <= x"00000000"; 
      when 4401 => DO <= x"00000000"; 
      when 4402 => DO <= x"00000000"; 
      when 4403 => DO <= x"00000000"; 
      when 4404 => DO <= x"00000000"; 
      when 4405 => DO <= x"00000000"; 
      when 4406 => DO <= x"00000000"; 
      when 4407 => DO <= x"00000000"; 
      when 4408 => DO <= x"00000000"; 
      when 4409 => DO <= x"00000000"; 
      when 4410 => DO <= x"00000000"; 
      when 4411 => DO <= x"00000000"; 
      when 4412 => DO <= x"00000000"; 
      when 4413 => DO <= x"00000000"; 
      when 4414 => DO <= x"00000000"; 
      when 4415 => DO <= x"00000000"; 
      when 4416 => DO <= x"00000000"; 
      when 4417 => DO <= x"00000000"; 
      when 4418 => DO <= x"00000000"; 
      when 4419 => DO <= x"00000000"; 
      when 4420 => DO <= x"00000000"; 
      when 4421 => DO <= x"00000000"; 
      when 4422 => DO <= x"00000000"; 
      when 4423 => DO <= x"00000000"; 
      when 4424 => DO <= x"00000000"; 
      when 4425 => DO <= x"00000000"; 
      when 4426 => DO <= x"00000000"; 
      when 4427 => DO <= x"00000000"; 
      when 4428 => DO <= x"00000000"; 
      when 4429 => DO <= x"00000000"; 
      when 4430 => DO <= x"00000000"; 
      when 4431 => DO <= x"00000000"; 
      when 4432 => DO <= x"00000000"; 
      when 4433 => DO <= x"00000000"; 
      when 4434 => DO <= x"00000000"; 
      when 4435 => DO <= x"00000000"; 
      when 4436 => DO <= x"00000000"; 
      when 4437 => DO <= x"00000000"; 
      when 4438 => DO <= x"00000000"; 
      when 4439 => DO <= x"00000000"; 
      when 4440 => DO <= x"00000000"; 
      when 4441 => DO <= x"00000000"; 
      when 4442 => DO <= x"00000000"; 
      when 4443 => DO <= x"00000000"; 
      when 4444 => DO <= x"00000000"; 
      when 4445 => DO <= x"00000000"; 
      when 4446 => DO <= x"00000000"; 
      when 4447 => DO <= x"00000000"; 
      when 4448 => DO <= x"00000000"; 
      when 4449 => DO <= x"00000000"; 
      when 4450 => DO <= x"00000000"; 
      when 4451 => DO <= x"00000000"; 
      when 4452 => DO <= x"00000000"; 
      when 4453 => DO <= x"00000000"; 
      when 4454 => DO <= x"00000000"; 
      when 4455 => DO <= x"00000000"; 
      when 4456 => DO <= x"00000000"; 
      when 4457 => DO <= x"00000000"; 
      when 4458 => DO <= x"00000000"; 
      when 4459 => DO <= x"00000000"; 
      when 4460 => DO <= x"00000000"; 
      when 4461 => DO <= x"00000000"; 
      when 4462 => DO <= x"00000000"; 
      when 4463 => DO <= x"00000000"; 
      when 4464 => DO <= x"00000000"; 
      when 4465 => DO <= x"00000000"; 
      when 4466 => DO <= x"00000000"; 
      when 4467 => DO <= x"00000000"; 
      when 4468 => DO <= x"00000000"; 
      when 4469 => DO <= x"00000000"; 
      when 4470 => DO <= x"00000000"; 
      when 4471 => DO <= x"00000000"; 
      when 4472 => DO <= x"00000000"; 
      when 4473 => DO <= x"00000000"; 
      when 4474 => DO <= x"00000000"; 
      when 4475 => DO <= x"00000000"; 
      when 4476 => DO <= x"00000000"; 
      when 4477 => DO <= x"00000000"; 
      when 4478 => DO <= x"00000000"; 
      when 4479 => DO <= x"00000000"; 
      when 4480 => DO <= x"00000000"; 
      when 4481 => DO <= x"00000000"; 
      when 4482 => DO <= x"00000000"; 
      when 4483 => DO <= x"00000000"; 
      when 4484 => DO <= x"00000000"; 
      when 4485 => DO <= x"00000000"; 
      when 4486 => DO <= x"00000000"; 
      when 4487 => DO <= x"00000000"; 
      when 4488 => DO <= x"00000000"; 
      when 4489 => DO <= x"00000000"; 
      when 4490 => DO <= x"00000000"; 
      when 4491 => DO <= x"00000000"; 
      when 4492 => DO <= x"00000000"; 
      when 4493 => DO <= x"00000000"; 
      when 4494 => DO <= x"00000000"; 
      when 4495 => DO <= x"00000000"; 
      when 4496 => DO <= x"00000000"; 
      when 4497 => DO <= x"00000000"; 
      when 4498 => DO <= x"00000000"; 
      when 4499 => DO <= x"00000000"; 
      when 4500 => DO <= x"00000000"; 
      when 4501 => DO <= x"00000000"; 
      when 4502 => DO <= x"00000000"; 
      when 4503 => DO <= x"00000000"; 
      when 4504 => DO <= x"00000000"; 
      when 4505 => DO <= x"00000000"; 
      when 4506 => DO <= x"00000000"; 
      when 4507 => DO <= x"00000000"; 
      when 4508 => DO <= x"00000000"; 
      when 4509 => DO <= x"00000000"; 
      when 4510 => DO <= x"00000000"; 
      when 4511 => DO <= x"00000000"; 
      when 4512 => DO <= x"00000000"; 
      when 4513 => DO <= x"00000000"; 
      when 4514 => DO <= x"00000000"; 
      when 4515 => DO <= x"00000000"; 
      when 4516 => DO <= x"00000000"; 
      when 4517 => DO <= x"00000000"; 
      when 4518 => DO <= x"00000000"; 
      when 4519 => DO <= x"00000000"; 
      when 4520 => DO <= x"00000000"; 
      when 4521 => DO <= x"00000000"; 
      when 4522 => DO <= x"00000000"; 
      when 4523 => DO <= x"00000000"; 
      when 4524 => DO <= x"00000000"; 
      when 4525 => DO <= x"00000000"; 
      when 4526 => DO <= x"00000000"; 
      when 4527 => DO <= x"00000000"; 
      when 4528 => DO <= x"00000000"; 
      when 4529 => DO <= x"00000000"; 
      when 4530 => DO <= x"00000000"; 
      when 4531 => DO <= x"00000000"; 
      when 4532 => DO <= x"00000000"; 
      when 4533 => DO <= x"00000000"; 
      when 4534 => DO <= x"00000000"; 
      when 4535 => DO <= x"00000000"; 
      when 4536 => DO <= x"00000000"; 
      when 4537 => DO <= x"00000000"; 
      when 4538 => DO <= x"00000000"; 
      when 4539 => DO <= x"00000000"; 
      when 4540 => DO <= x"00000000"; 
      when 4541 => DO <= x"00000000"; 
      when 4542 => DO <= x"00000000"; 
      when 4543 => DO <= x"00000000"; 
      when 4544 => DO <= x"00000000"; 
      when 4545 => DO <= x"00000000"; 
      when 4546 => DO <= x"00000000"; 
      when 4547 => DO <= x"00000000"; 
      when 4548 => DO <= x"00000000"; 
      when 4549 => DO <= x"00000000"; 
      when 4550 => DO <= x"00000000"; 
      when 4551 => DO <= x"00000000"; 
      when 4552 => DO <= x"00000000"; 
      when 4553 => DO <= x"00000000"; 
      when 4554 => DO <= x"00000000"; 
      when 4555 => DO <= x"00000000"; 
      when 4556 => DO <= x"00000000"; 
      when 4557 => DO <= x"00000000"; 
      when 4558 => DO <= x"00000000"; 
      when 4559 => DO <= x"00000000"; 
      when 4560 => DO <= x"00000000"; 
      when 4561 => DO <= x"00000000"; 
      when 4562 => DO <= x"00000000"; 
      when 4563 => DO <= x"00000000"; 
      when 4564 => DO <= x"00000000"; 
      when 4565 => DO <= x"00000000"; 
      when 4566 => DO <= x"00000000"; 
      when 4567 => DO <= x"00000000"; 
      when 4568 => DO <= x"00000000"; 
      when 4569 => DO <= x"00000000"; 
      when 4570 => DO <= x"00000000"; 
      when 4571 => DO <= x"00000000"; 
      when 4572 => DO <= x"00000000"; 
      when 4573 => DO <= x"00000000"; 
      when 4574 => DO <= x"00000000"; 
      when 4575 => DO <= x"00000000"; 
      when 4576 => DO <= x"00000000"; 
      when 4577 => DO <= x"00000000"; 
      when 4578 => DO <= x"00000000"; 
      when 4579 => DO <= x"00000000"; 
      when 4580 => DO <= x"00000000"; 
      when 4581 => DO <= x"00000000"; 
      when 4582 => DO <= x"00000000"; 
      when 4583 => DO <= x"00000000"; 
      when 4584 => DO <= x"00000000"; 
      when 4585 => DO <= x"00000000"; 
      when 4586 => DO <= x"00000000"; 
      when 4587 => DO <= x"00000000"; 
      when 4588 => DO <= x"00000000"; 
      when 4589 => DO <= x"00000000"; 
      when 4590 => DO <= x"00000000"; 
      when 4591 => DO <= x"00000000"; 
      when 4592 => DO <= x"00000000"; 
      when 4593 => DO <= x"00000000"; 
      when 4594 => DO <= x"00000000"; 
      when 4595 => DO <= x"00000000"; 
      when 4596 => DO <= x"00000000"; 
      when 4597 => DO <= x"00000000"; 
      when 4598 => DO <= x"00000000"; 
      when 4599 => DO <= x"00000000"; 
      when 4600 => DO <= x"00000000"; 
      when 4601 => DO <= x"00000000"; 
      when 4602 => DO <= x"00000000"; 
      when 4603 => DO <= x"00000000"; 
      when 4604 => DO <= x"00000000"; 
      when 4605 => DO <= x"00000000"; 
      when 4606 => DO <= x"00000000"; 
      when 4607 => DO <= x"00000000"; 
      when 4608 => DO <= x"00000000"; 
      when 4609 => DO <= x"00000000"; 
      when 4610 => DO <= x"00000000"; 
      when 4611 => DO <= x"00000000"; 
      when 4612 => DO <= x"00000000"; 
      when 4613 => DO <= x"00000000"; 
      when 4614 => DO <= x"00000000"; 
      when 4615 => DO <= x"00000000"; 
      when 4616 => DO <= x"00000000"; 
      when 4617 => DO <= x"00000000"; 
      when 4618 => DO <= x"00000000"; 
      when 4619 => DO <= x"00000000"; 
      when 4620 => DO <= x"00000000"; 
      when 4621 => DO <= x"00000000"; 
      when 4622 => DO <= x"00000000"; 
      when 4623 => DO <= x"00000000"; 
      when 4624 => DO <= x"00000000"; 
      when 4625 => DO <= x"00000000"; 
      when 4626 => DO <= x"00000000"; 
      when 4627 => DO <= x"00000000"; 
      when 4628 => DO <= x"00000000"; 
      when 4629 => DO <= x"00000000"; 
      when 4630 => DO <= x"00000000"; 
      when 4631 => DO <= x"00000000"; 
      when 4632 => DO <= x"00000000"; 
      when 4633 => DO <= x"00000000"; 
      when 4634 => DO <= x"00000000"; 
      when 4635 => DO <= x"00000000"; 
      when 4636 => DO <= x"00000000"; 
      when 4637 => DO <= x"00000000"; 
      when 4638 => DO <= x"00000000"; 
      when 4639 => DO <= x"00000000"; 
      when 4640 => DO <= x"00000000"; 
      when 4641 => DO <= x"00000000"; 
      when 4642 => DO <= x"00000000"; 
      when 4643 => DO <= x"00000000"; 
      when 4644 => DO <= x"00000000"; 
      when 4645 => DO <= x"00000000"; 
      when 4646 => DO <= x"00000000"; 
      when 4647 => DO <= x"00000000"; 
      when 4648 => DO <= x"00000000"; 
      when 4649 => DO <= x"00000000"; 
      when 4650 => DO <= x"00000000"; 
      when 4651 => DO <= x"00000000"; 
      when 4652 => DO <= x"00000000"; 
      when 4653 => DO <= x"00000000"; 
      when 4654 => DO <= x"00000000"; 
      when 4655 => DO <= x"00000000"; 
      when 4656 => DO <= x"00000000"; 
      when 4657 => DO <= x"00000000"; 
      when 4658 => DO <= x"00000000"; 
      when 4659 => DO <= x"00000000"; 
      when 4660 => DO <= x"00000000"; 
      when 4661 => DO <= x"00000000"; 
      when 4662 => DO <= x"00000000"; 
      when 4663 => DO <= x"00000000"; 
      when 4664 => DO <= x"00000000"; 
      when 4665 => DO <= x"00000000"; 
      when 4666 => DO <= x"00000000"; 
      when 4667 => DO <= x"00000000"; 
      when 4668 => DO <= x"00000000"; 
      when 4669 => DO <= x"00000000"; 
      when 4670 => DO <= x"00000000"; 
      when 4671 => DO <= x"00000000"; 
      when 4672 => DO <= x"00000000"; 
      when 4673 => DO <= x"00000000"; 
      when 4674 => DO <= x"00000000"; 
      when 4675 => DO <= x"00000000"; 
      when 4676 => DO <= x"00000000"; 
      when 4677 => DO <= x"00000000"; 
      when 4678 => DO <= x"00000000"; 
      when 4679 => DO <= x"00000000"; 
      when 4680 => DO <= x"00000000"; 
      when 4681 => DO <= x"00000000"; 
      when 4682 => DO <= x"00000000"; 
      when 4683 => DO <= x"00000000"; 
      when 4684 => DO <= x"00000000"; 
      when 4685 => DO <= x"00000000"; 
      when 4686 => DO <= x"00000000"; 
      when 4687 => DO <= x"00000000"; 
      when 4688 => DO <= x"00000000"; 
      when 4689 => DO <= x"00000000"; 
      when 4690 => DO <= x"00000000"; 
      when 4691 => DO <= x"00000000"; 
      when 4692 => DO <= x"00000000"; 
      when 4693 => DO <= x"00000000"; 
      when 4694 => DO <= x"00000000"; 
      when 4695 => DO <= x"00000000"; 
      when 4696 => DO <= x"00000000"; 
      when 4697 => DO <= x"00000000"; 
      when 4698 => DO <= x"00000000"; 
      when 4699 => DO <= x"00000000"; 
      when 4700 => DO <= x"00000000"; 
      when 4701 => DO <= x"00000000"; 
      when 4702 => DO <= x"00000000"; 
      when 4703 => DO <= x"00000000"; 
      when 4704 => DO <= x"00000000"; 
      when 4705 => DO <= x"00000000"; 
      when 4706 => DO <= x"00000000"; 
      when 4707 => DO <= x"00000000"; 
      when 4708 => DO <= x"00000000"; 
      when 4709 => DO <= x"00000000"; 
      when 4710 => DO <= x"00000000"; 
      when 4711 => DO <= x"00000000"; 
      when 4712 => DO <= x"00000000"; 
      when 4713 => DO <= x"00000000"; 
      when 4714 => DO <= x"00000000"; 
      when 4715 => DO <= x"00000000"; 
      when 4716 => DO <= x"00000000"; 
      when 4717 => DO <= x"00000000"; 
      when 4718 => DO <= x"00000000"; 
      when 4719 => DO <= x"00000000"; 
      when 4720 => DO <= x"00000000"; 
      when 4721 => DO <= x"00000000"; 
      when 4722 => DO <= x"00000000"; 
      when 4723 => DO <= x"00000000"; 
      when 4724 => DO <= x"00000000"; 
      when 4725 => DO <= x"00000000"; 
      when 4726 => DO <= x"00000000"; 
      when 4727 => DO <= x"00000000"; 
      when 4728 => DO <= x"00000000"; 
      when 4729 => DO <= x"00000000"; 
      when 4730 => DO <= x"00000000"; 
      when 4731 => DO <= x"00000000"; 
      when 4732 => DO <= x"00000000"; 
      when 4733 => DO <= x"00000000"; 
      when 4734 => DO <= x"00000000"; 
      when 4735 => DO <= x"00000000"; 
      when 4736 => DO <= x"00000000"; 
      when 4737 => DO <= x"00000000"; 
      when 4738 => DO <= x"00000000"; 
      when 4739 => DO <= x"00000000"; 
      when 4740 => DO <= x"00000000"; 
      when 4741 => DO <= x"00000000"; 
      when 4742 => DO <= x"00000000"; 
      when 4743 => DO <= x"00000000"; 
      when 4744 => DO <= x"00000000"; 
      when 4745 => DO <= x"00000000"; 
      when 4746 => DO <= x"00000000"; 
      when 4747 => DO <= x"00000000"; 
      when 4748 => DO <= x"00000000"; 
      when 4749 => DO <= x"00000000"; 
      when 4750 => DO <= x"00000000"; 
      when 4751 => DO <= x"00000000"; 
      when 4752 => DO <= x"00000000"; 
      when 4753 => DO <= x"00000000"; 
      when 4754 => DO <= x"00000000"; 
      when 4755 => DO <= x"00000000"; 
      when 4756 => DO <= x"00000000"; 
      when 4757 => DO <= x"00000000"; 
      when 4758 => DO <= x"00000000"; 
      when 4759 => DO <= x"00000000"; 
      when 4760 => DO <= x"00000000"; 
      when 4761 => DO <= x"00000000"; 
      when 4762 => DO <= x"00000000"; 
      when 4763 => DO <= x"00000000"; 
      when 4764 => DO <= x"00000000"; 
      when 4765 => DO <= x"00000000"; 
      when 4766 => DO <= x"00000000"; 
      when 4767 => DO <= x"00000000"; 
      when 4768 => DO <= x"00000000"; 
      when 4769 => DO <= x"00000000"; 
      when 4770 => DO <= x"00000000"; 
      when 4771 => DO <= x"00000000"; 
      when 4772 => DO <= x"00000000"; 
      when 4773 => DO <= x"00000000"; 
      when 4774 => DO <= x"00000000"; 
      when 4775 => DO <= x"00000000"; 
      when 4776 => DO <= x"00000000"; 
      when 4777 => DO <= x"00000000"; 
      when 4778 => DO <= x"00000000"; 
      when 4779 => DO <= x"00000000"; 
      when 4780 => DO <= x"00000000"; 
      when 4781 => DO <= x"00000000"; 
      when 4782 => DO <= x"00000000"; 
      when 4783 => DO <= x"00000000"; 
      when 4784 => DO <= x"00000000"; 
      when 4785 => DO <= x"00000000"; 
      when 4786 => DO <= x"00000000"; 
      when 4787 => DO <= x"00000000"; 
      when 4788 => DO <= x"00000000"; 
      when 4789 => DO <= x"00000000"; 
      when 4790 => DO <= x"00000000"; 
      when 4791 => DO <= x"00000000"; 
      when 4792 => DO <= x"00000000"; 
      when 4793 => DO <= x"00000000"; 
      when 4794 => DO <= x"00000000"; 
      when 4795 => DO <= x"00000000"; 
      when 4796 => DO <= x"00000000"; 
      when 4797 => DO <= x"00000000"; 
      when 4798 => DO <= x"00000000"; 
      when 4799 => DO <= x"00000000"; 
      when 4800 => DO <= x"00000000"; 
      when 4801 => DO <= x"00000000"; 
      when 4802 => DO <= x"00000000"; 
      when 4803 => DO <= x"00000000"; 
      when 4804 => DO <= x"00000000"; 
      when 4805 => DO <= x"00000000"; 
      when 4806 => DO <= x"00000000"; 
      when 4807 => DO <= x"00000000"; 
      when 4808 => DO <= x"00000000"; 
      when 4809 => DO <= x"00000000"; 
      when 4810 => DO <= x"00000000"; 
      when 4811 => DO <= x"00000000"; 
      when 4812 => DO <= x"00000000"; 
      when 4813 => DO <= x"00000000"; 
      when 4814 => DO <= x"00000000"; 
      when 4815 => DO <= x"00000000"; 
      when 4816 => DO <= x"00000000"; 
      when 4817 => DO <= x"00000000"; 
      when 4818 => DO <= x"00000000"; 
      when 4819 => DO <= x"00000000"; 
      when 4820 => DO <= x"00000000"; 
      when 4821 => DO <= x"00000000"; 
      when 4822 => DO <= x"00000000"; 
      when 4823 => DO <= x"00000000"; 
      when 4824 => DO <= x"00000000"; 
      when 4825 => DO <= x"00000000"; 
      when 4826 => DO <= x"00000000"; 
      when 4827 => DO <= x"00000000"; 
      when 4828 => DO <= x"00000000"; 
      when 4829 => DO <= x"00000000"; 
      when 4830 => DO <= x"00000000"; 
      when 4831 => DO <= x"00000000"; 
      when 4832 => DO <= x"00000000"; 
      when 4833 => DO <= x"00000000"; 
      when 4834 => DO <= x"00000000"; 
      when 4835 => DO <= x"00000000"; 
      when 4836 => DO <= x"00000000"; 
      when 4837 => DO <= x"00000000"; 
      when 4838 => DO <= x"00000000"; 
      when 4839 => DO <= x"00000000"; 
      when 4840 => DO <= x"00000000"; 
      when 4841 => DO <= x"00000000"; 
      when 4842 => DO <= x"00000000"; 
      when 4843 => DO <= x"00000000"; 
      when 4844 => DO <= x"00000000"; 
      when 4845 => DO <= x"00000000"; 
      when 4846 => DO <= x"00000000"; 
      when 4847 => DO <= x"00000000"; 
      when 4848 => DO <= x"00000000"; 
      when 4849 => DO <= x"00000000"; 
      when 4850 => DO <= x"00000000"; 
      when 4851 => DO <= x"00000000"; 
      when 4852 => DO <= x"00000000"; 
      when 4853 => DO <= x"00000000"; 
      when 4854 => DO <= x"00000000"; 
      when 4855 => DO <= x"00000000"; 
      when 4856 => DO <= x"00000000"; 
      when 4857 => DO <= x"00000000"; 
      when 4858 => DO <= x"00000000"; 
      when 4859 => DO <= x"00000000"; 
      when 4860 => DO <= x"00000000"; 
      when 4861 => DO <= x"00000000"; 
      when 4862 => DO <= x"00000000"; 
      when 4863 => DO <= x"00000000"; 
      when 4864 => DO <= x"00000000"; 
      when 4865 => DO <= x"00000000"; 
      when 4866 => DO <= x"00000000"; 
      when 4867 => DO <= x"00000000"; 
      when 4868 => DO <= x"00000000"; 
      when 4869 => DO <= x"00000000"; 
      when 4870 => DO <= x"00000000"; 
      when 4871 => DO <= x"00000000"; 
      when 4872 => DO <= x"00000000"; 
      when 4873 => DO <= x"00000000"; 
      when 4874 => DO <= x"00000000"; 
      when 4875 => DO <= x"00000000"; 
      when 4876 => DO <= x"00000000"; 
      when 4877 => DO <= x"00000000"; 
      when 4878 => DO <= x"00000000"; 
      when 4879 => DO <= x"00000000"; 
      when 4880 => DO <= x"00000000"; 
      when 4881 => DO <= x"00000000"; 
      when 4882 => DO <= x"00000000"; 
      when 4883 => DO <= x"00000000"; 
      when 4884 => DO <= x"00000000"; 
      when 4885 => DO <= x"00000000"; 
      when 4886 => DO <= x"00000000"; 
      when 4887 => DO <= x"00000000"; 
      when 4888 => DO <= x"00000000"; 
      when 4889 => DO <= x"00000000"; 
      when 4890 => DO <= x"00000000"; 
      when 4891 => DO <= x"00000000"; 
      when 4892 => DO <= x"00000000"; 
      when 4893 => DO <= x"00000000"; 
      when 4894 => DO <= x"00000000"; 
      when 4895 => DO <= x"00000000"; 
      when 4896 => DO <= x"00000000"; 
      when 4897 => DO <= x"00000000"; 
      when 4898 => DO <= x"00000000"; 
      when 4899 => DO <= x"00000000"; 
      when 4900 => DO <= x"00000000"; 
      when 4901 => DO <= x"00000000"; 
      when 4902 => DO <= x"00000000"; 
      when 4903 => DO <= x"00000000"; 
      when 4904 => DO <= x"00000000"; 
      when 4905 => DO <= x"00000000"; 
      when 4906 => DO <= x"00000000"; 
      when 4907 => DO <= x"00000000"; 
      when 4908 => DO <= x"00000000"; 
      when 4909 => DO <= x"00000000"; 
      when 4910 => DO <= x"00000000"; 
      when 4911 => DO <= x"00000000"; 
      when 4912 => DO <= x"00000000"; 
      when 4913 => DO <= x"00000000"; 
      when 4914 => DO <= x"00000000"; 
      when 4915 => DO <= x"00000000"; 
      when 4916 => DO <= x"00000000"; 
      when 4917 => DO <= x"00000000"; 
      when 4918 => DO <= x"00000000"; 
      when 4919 => DO <= x"00000000"; 
      when 4920 => DO <= x"00000000"; 
      when 4921 => DO <= x"00000000"; 
      when 4922 => DO <= x"00000000"; 
      when 4923 => DO <= x"00000000"; 
      when 4924 => DO <= x"00000000"; 
      when 4925 => DO <= x"00000000"; 
      when 4926 => DO <= x"00000000"; 
      when 4927 => DO <= x"00000000"; 
      when 4928 => DO <= x"00000000"; 
      when 4929 => DO <= x"00000000"; 
      when 4930 => DO <= x"00000000"; 
      when 4931 => DO <= x"00000000"; 
      when 4932 => DO <= x"00000000"; 
      when 4933 => DO <= x"00000000"; 
      when 4934 => DO <= x"00000000"; 
      when 4935 => DO <= x"00000000"; 
      when 4936 => DO <= x"00000000"; 
      when 4937 => DO <= x"00000000"; 
      when 4938 => DO <= x"00000000"; 
      when 4939 => DO <= x"00000000"; 
      when 4940 => DO <= x"00000000"; 
      when 4941 => DO <= x"00000000"; 
      when 4942 => DO <= x"00000000"; 
      when 4943 => DO <= x"00000000"; 
      when 4944 => DO <= x"00000000"; 
      when 4945 => DO <= x"00000000"; 
      when 4946 => DO <= x"00000000"; 
      when 4947 => DO <= x"00000000"; 
      when 4948 => DO <= x"00000000"; 
      when 4949 => DO <= x"00000000"; 
      when 4950 => DO <= x"00000000"; 
      when 4951 => DO <= x"00000000"; 
      when 4952 => DO <= x"00000000"; 
      when 4953 => DO <= x"00000000"; 
      when 4954 => DO <= x"00000000"; 
      when 4955 => DO <= x"00000000"; 
      when 4956 => DO <= x"00000000"; 
      when 4957 => DO <= x"00000000"; 
      when 4958 => DO <= x"00000000"; 
      when 4959 => DO <= x"00000000"; 
      when 4960 => DO <= x"00000000"; 
      when 4961 => DO <= x"00000000"; 
      when 4962 => DO <= x"00000000"; 
      when 4963 => DO <= x"00000000"; 
      when 4964 => DO <= x"00000000"; 
      when 4965 => DO <= x"00000000"; 
      when 4966 => DO <= x"00000000"; 
      when 4967 => DO <= x"00000000"; 
      when 4968 => DO <= x"00000000"; 
      when 4969 => DO <= x"00000000"; 
      when 4970 => DO <= x"00000000"; 
      when 4971 => DO <= x"00000000"; 
      when 4972 => DO <= x"00000000"; 
      when 4973 => DO <= x"00000000"; 
      when 4974 => DO <= x"00000000"; 
      when 4975 => DO <= x"00000000"; 
      when 4976 => DO <= x"00000000"; 
      when 4977 => DO <= x"00000000"; 
      when 4978 => DO <= x"00000000"; 
      when 4979 => DO <= x"00000000"; 
      when 4980 => DO <= x"00000000"; 
      when 4981 => DO <= x"00000000"; 
      when 4982 => DO <= x"00000000"; 
      when 4983 => DO <= x"00000000"; 
      when 4984 => DO <= x"00000000"; 
      when 4985 => DO <= x"00000000"; 
      when 4986 => DO <= x"00000000"; 
      when 4987 => DO <= x"00000000"; 
      when 4988 => DO <= x"00000000"; 
      when 4989 => DO <= x"00000000"; 
      when 4990 => DO <= x"00000000"; 
      when 4991 => DO <= x"00000000"; 
      when 4992 => DO <= x"00000000"; 
      when 4993 => DO <= x"00000000"; 
      when 4994 => DO <= x"00000000"; 
      when 4995 => DO <= x"00000000"; 
      when 4996 => DO <= x"00000000"; 
      when 4997 => DO <= x"00000000"; 
      when 4998 => DO <= x"00000000"; 
      when 4999 => DO <= x"00000000"; 
      when 5000 => DO <= x"00000000"; 
      when 5001 => DO <= x"00000000"; 
      when 5002 => DO <= x"00000000"; 
      when 5003 => DO <= x"00000000"; 
      when 5004 => DO <= x"00000000"; 
      when 5005 => DO <= x"00000000"; 
      when 5006 => DO <= x"00000000"; 
      when 5007 => DO <= x"00000000"; 
      when 5008 => DO <= x"00000000"; 
      when 5009 => DO <= x"00000000"; 
      when 5010 => DO <= x"00000000"; 
      when 5011 => DO <= x"00000000"; 
      when 5012 => DO <= x"00000000"; 
      when 5013 => DO <= x"00000000"; 
      when 5014 => DO <= x"00000000"; 
      when 5015 => DO <= x"00000000"; 
      when 5016 => DO <= x"00000000"; 
      when 5017 => DO <= x"00000000"; 
      when 5018 => DO <= x"00000000"; 
      when 5019 => DO <= x"00000000"; 
      when 5020 => DO <= x"00000000"; 
      when 5021 => DO <= x"00000000"; 
      when 5022 => DO <= x"00000000"; 
      when 5023 => DO <= x"00000000"; 
      when 5024 => DO <= x"00000000"; 
      when 5025 => DO <= x"00000000"; 
      when 5026 => DO <= x"00000000"; 
      when 5027 => DO <= x"00000000"; 
      when 5028 => DO <= x"00000000"; 
      when 5029 => DO <= x"00000000"; 
      when 5030 => DO <= x"00000000"; 
      when 5031 => DO <= x"00000000"; 
      when 5032 => DO <= x"00000000"; 
      when 5033 => DO <= x"00000000"; 
      when 5034 => DO <= x"00000000"; 
      when 5035 => DO <= x"00000000"; 
      when 5036 => DO <= x"00000000"; 
      when 5037 => DO <= x"00000000"; 
      when 5038 => DO <= x"00000000"; 
      when 5039 => DO <= x"00000000"; 
      when 5040 => DO <= x"00000000"; 
      when 5041 => DO <= x"00000000"; 
      when 5042 => DO <= x"00000000"; 
      when 5043 => DO <= x"00000000"; 
      when 5044 => DO <= x"00000000"; 
      when 5045 => DO <= x"00000000"; 
      when 5046 => DO <= x"00000000"; 
      when 5047 => DO <= x"00000000"; 
      when 5048 => DO <= x"00000000"; 
      when 5049 => DO <= x"00000000"; 
      when 5050 => DO <= x"00000000"; 
      when 5051 => DO <= x"00000000"; 
      when 5052 => DO <= x"00000000"; 
      when 5053 => DO <= x"00000000"; 
      when 5054 => DO <= x"00000000"; 
      when 5055 => DO <= x"00000000"; 
      when 5056 => DO <= x"00000000"; 
      when 5057 => DO <= x"00000000"; 
      when 5058 => DO <= x"00000000"; 
      when 5059 => DO <= x"00000000"; 
      when 5060 => DO <= x"00000000"; 
      when 5061 => DO <= x"00000000"; 
      when 5062 => DO <= x"00000000"; 
      when 5063 => DO <= x"00000000"; 
      when 5064 => DO <= x"00000000"; 
      when 5065 => DO <= x"00000000"; 
      when 5066 => DO <= x"00000000"; 
      when 5067 => DO <= x"00000000"; 
      when 5068 => DO <= x"00000000"; 
      when 5069 => DO <= x"00000000"; 
      when 5070 => DO <= x"00000000"; 
      when 5071 => DO <= x"00000000"; 
      when 5072 => DO <= x"00000000"; 
      when 5073 => DO <= x"00000000"; 
      when 5074 => DO <= x"00000000"; 
      when 5075 => DO <= x"00000000"; 
      when 5076 => DO <= x"00000000"; 
      when 5077 => DO <= x"00000000"; 
      when 5078 => DO <= x"00000000"; 
      when 5079 => DO <= x"00000000"; 
      when 5080 => DO <= x"00000000"; 
      when 5081 => DO <= x"00000000"; 
      when 5082 => DO <= x"00000000"; 
      when 5083 => DO <= x"00000000"; 
      when 5084 => DO <= x"00000000"; 
      when 5085 => DO <= x"00000000"; 
      when 5086 => DO <= x"00000000"; 
      when 5087 => DO <= x"00000000"; 
      when 5088 => DO <= x"00000000"; 
      when 5089 => DO <= x"00000000"; 
      when 5090 => DO <= x"00000000"; 
      when 5091 => DO <= x"00000000"; 
      when 5092 => DO <= x"00000000"; 
      when 5093 => DO <= x"00000000"; 
      when 5094 => DO <= x"00000000"; 
      when 5095 => DO <= x"00000000"; 
      when 5096 => DO <= x"00000000"; 
      when 5097 => DO <= x"00000000"; 
      when 5098 => DO <= x"00000000"; 
      when 5099 => DO <= x"00000000"; 
      when 5100 => DO <= x"00000000"; 
      when 5101 => DO <= x"00000000"; 
      when 5102 => DO <= x"00000000"; 
      when 5103 => DO <= x"00000000"; 
      when 5104 => DO <= x"00000000"; 
      when 5105 => DO <= x"00000000"; 
      when 5106 => DO <= x"00000000"; 
      when 5107 => DO <= x"00000000"; 
      when 5108 => DO <= x"00000000"; 
      when 5109 => DO <= x"00000000"; 
      when 5110 => DO <= x"00000000"; 
      when 5111 => DO <= x"00000000"; 
      when 5112 => DO <= x"00000000"; 
      when 5113 => DO <= x"00000000"; 
      when 5114 => DO <= x"00000000"; 
      when 5115 => DO <= x"00000000"; 
      when 5116 => DO <= x"00000000"; 
      when 5117 => DO <= x"00000000"; 
      when 5118 => DO <= x"00000000"; 
      when 5119 => DO <= x"00000000"; 
      when 5120 => DO <= x"00000000"; 
      when 5121 => DO <= x"00000000"; 
      when 5122 => DO <= x"00000000"; 
      when 5123 => DO <= x"00000000"; 
      when 5124 => DO <= x"00000000"; 
      when 5125 => DO <= x"00000000"; 
      when 5126 => DO <= x"00000000"; 
      when 5127 => DO <= x"00000000"; 
      when 5128 => DO <= x"00000000"; 
      when 5129 => DO <= x"00000000"; 
      when 5130 => DO <= x"00000000"; 
      when 5131 => DO <= x"00000000"; 
      when 5132 => DO <= x"00000000"; 
      when 5133 => DO <= x"00000000"; 
      when 5134 => DO <= x"00000000"; 
      when 5135 => DO <= x"00000000"; 
      when 5136 => DO <= x"00000000"; 
      when 5137 => DO <= x"00000000"; 
      when 5138 => DO <= x"00000000"; 
      when 5139 => DO <= x"00000000"; 
      when 5140 => DO <= x"00000000"; 
      when 5141 => DO <= x"00000000"; 
      when 5142 => DO <= x"00000000"; 
      when 5143 => DO <= x"00000000"; 
      when 5144 => DO <= x"00000000"; 
      when 5145 => DO <= x"00000000"; 
      when 5146 => DO <= x"00000000"; 
      when 5147 => DO <= x"00000000"; 
      when 5148 => DO <= x"00000000"; 
      when 5149 => DO <= x"00000000"; 
      when 5150 => DO <= x"00000000"; 
      when 5151 => DO <= x"00000000"; 
      when 5152 => DO <= x"00000000"; 
      when 5153 => DO <= x"00000000"; 
      when 5154 => DO <= x"00000000"; 
      when 5155 => DO <= x"00000000"; 
      when 5156 => DO <= x"00000000"; 
      when 5157 => DO <= x"00000000"; 
      when 5158 => DO <= x"00000000"; 
      when 5159 => DO <= x"00000000"; 
      when 5160 => DO <= x"00000000"; 
      when 5161 => DO <= x"00000000"; 
      when 5162 => DO <= x"00000000"; 
      when 5163 => DO <= x"00000000"; 
      when 5164 => DO <= x"00000000"; 
      when 5165 => DO <= x"00000000"; 
      when 5166 => DO <= x"00000000"; 
      when 5167 => DO <= x"00000000"; 
      when 5168 => DO <= x"00000000"; 
      when 5169 => DO <= x"00000000"; 
      when 5170 => DO <= x"00000000"; 
      when 5171 => DO <= x"00000000"; 
      when 5172 => DO <= x"00000000"; 
      when 5173 => DO <= x"00000000"; 
      when 5174 => DO <= x"00000000"; 
      when 5175 => DO <= x"00000000"; 
      when 5176 => DO <= x"00000000"; 
      when 5177 => DO <= x"00000000"; 
      when 5178 => DO <= x"00000000"; 
      when 5179 => DO <= x"00000000"; 
      when 5180 => DO <= x"00000000"; 
      when 5181 => DO <= x"00000000"; 
      when 5182 => DO <= x"00000000"; 
      when 5183 => DO <= x"00000000"; 
      when 5184 => DO <= x"00000000"; 
      when 5185 => DO <= x"00000000"; 
      when 5186 => DO <= x"00000000"; 
      when 5187 => DO <= x"00000000"; 
      when 5188 => DO <= x"00000000"; 
      when 5189 => DO <= x"00000000"; 
      when 5190 => DO <= x"00000000"; 
      when 5191 => DO <= x"00000000"; 
      when 5192 => DO <= x"00000000"; 
      when 5193 => DO <= x"00000000"; 
      when 5194 => DO <= x"00000000"; 
      when 5195 => DO <= x"00000000"; 
      when 5196 => DO <= x"00000000"; 
      when 5197 => DO <= x"00000000"; 
      when 5198 => DO <= x"00000000"; 
      when 5199 => DO <= x"00000000"; 
      when 5200 => DO <= x"00000000"; 
      when 5201 => DO <= x"00000000"; 
      when 5202 => DO <= x"00000000"; 
      when 5203 => DO <= x"00000000"; 
      when 5204 => DO <= x"00000000"; 
      when 5205 => DO <= x"00000000"; 
      when 5206 => DO <= x"00000000"; 
      when 5207 => DO <= x"00000000"; 
      when 5208 => DO <= x"00000000"; 
      when 5209 => DO <= x"00000000"; 
      when 5210 => DO <= x"00000000"; 
      when 5211 => DO <= x"00000000"; 
      when 5212 => DO <= x"00000000"; 
      when 5213 => DO <= x"00000000"; 
      when 5214 => DO <= x"00000000"; 
      when 5215 => DO <= x"00000000"; 
      when 5216 => DO <= x"00000000"; 
      when 5217 => DO <= x"00000000"; 
      when 5218 => DO <= x"00000000"; 
      when 5219 => DO <= x"00000000"; 
      when 5220 => DO <= x"00000000"; 
      when 5221 => DO <= x"00000000"; 
      when 5222 => DO <= x"00000000"; 
      when 5223 => DO <= x"00000000"; 
      when 5224 => DO <= x"00000000"; 
      when 5225 => DO <= x"00000000"; 
      when 5226 => DO <= x"00000000"; 
      when 5227 => DO <= x"00000000"; 
      when 5228 => DO <= x"00000000"; 
      when 5229 => DO <= x"00000000"; 
      when 5230 => DO <= x"00000000"; 
      when 5231 => DO <= x"00000000"; 
      when 5232 => DO <= x"00000000"; 
      when 5233 => DO <= x"00000000"; 
      when 5234 => DO <= x"00000000"; 
      when 5235 => DO <= x"00000000"; 
      when 5236 => DO <= x"00000000"; 
      when 5237 => DO <= x"00000000"; 
      when 5238 => DO <= x"00000000"; 
      when 5239 => DO <= x"00000000"; 
      when 5240 => DO <= x"00000000"; 
      when 5241 => DO <= x"00000000"; 
      when 5242 => DO <= x"00000000"; 
      when 5243 => DO <= x"00000000"; 
      when 5244 => DO <= x"00000000"; 
      when 5245 => DO <= x"00000000"; 
      when 5246 => DO <= x"00000000"; 
      when 5247 => DO <= x"00000000"; 
      when 5248 => DO <= x"00000000"; 
      when 5249 => DO <= x"00000000"; 
      when 5250 => DO <= x"00000000"; 
      when 5251 => DO <= x"00000000"; 
      when 5252 => DO <= x"00000000"; 
      when 5253 => DO <= x"00000000"; 
      when 5254 => DO <= x"00000000"; 
      when 5255 => DO <= x"00000000"; 
      when 5256 => DO <= x"00000000"; 
      when 5257 => DO <= x"00000000"; 
      when 5258 => DO <= x"00000000"; 
      when 5259 => DO <= x"00000000"; 
      when 5260 => DO <= x"00000000"; 
      when 5261 => DO <= x"00000000"; 
      when 5262 => DO <= x"00000000"; 
      when 5263 => DO <= x"00000000"; 
      when 5264 => DO <= x"00000000"; 
      when 5265 => DO <= x"00000000"; 
      when 5266 => DO <= x"00000000"; 
      when 5267 => DO <= x"00000000"; 
      when 5268 => DO <= x"00000000"; 
      when 5269 => DO <= x"00000000"; 
      when 5270 => DO <= x"00000000"; 
      when 5271 => DO <= x"00000000"; 
      when 5272 => DO <= x"00000000"; 
      when 5273 => DO <= x"00000000"; 
      when 5274 => DO <= x"00000000"; 
      when 5275 => DO <= x"00000000"; 
      when 5276 => DO <= x"00000000"; 
      when 5277 => DO <= x"00000000"; 
      when 5278 => DO <= x"00000000"; 
      when 5279 => DO <= x"00000000"; 
      when 5280 => DO <= x"00000000"; 
      when 5281 => DO <= x"00000000"; 
      when 5282 => DO <= x"00000000"; 
      when 5283 => DO <= x"00000000"; 
      when 5284 => DO <= x"00000000"; 
      when 5285 => DO <= x"00000000"; 
      when 5286 => DO <= x"00000000"; 
      when 5287 => DO <= x"00000000"; 
      when 5288 => DO <= x"00000000"; 
      when 5289 => DO <= x"00000000"; 
      when 5290 => DO <= x"00000000"; 
      when 5291 => DO <= x"00000000"; 
      when 5292 => DO <= x"00000000"; 
      when 5293 => DO <= x"00000000"; 
      when 5294 => DO <= x"00000000"; 
      when 5295 => DO <= x"00000000"; 
      when 5296 => DO <= x"00000000"; 
      when 5297 => DO <= x"00000000"; 
      when 5298 => DO <= x"00000000"; 
      when 5299 => DO <= x"00000000"; 
      when 5300 => DO <= x"00000000"; 
      when 5301 => DO <= x"00000000"; 
      when 5302 => DO <= x"00000000"; 
      when 5303 => DO <= x"00000000"; 
      when 5304 => DO <= x"00000000"; 
      when 5305 => DO <= x"00000000"; 
      when 5306 => DO <= x"00000000"; 
      when 5307 => DO <= x"00000000"; 
      when 5308 => DO <= x"00000000"; 
      when 5309 => DO <= x"00000000"; 
      when 5310 => DO <= x"00000000"; 
      when 5311 => DO <= x"00000000"; 
      when 5312 => DO <= x"00000000"; 
      when 5313 => DO <= x"00000000"; 
      when 5314 => DO <= x"00000000"; 
      when 5315 => DO <= x"00000000"; 
      when 5316 => DO <= x"00000000"; 
      when 5317 => DO <= x"00000000"; 
      when 5318 => DO <= x"00000000"; 
      when 5319 => DO <= x"00000000"; 
      when 5320 => DO <= x"00000000"; 
      when 5321 => DO <= x"00000000"; 
      when 5322 => DO <= x"00000000"; 
      when 5323 => DO <= x"00000000"; 
      when 5324 => DO <= x"00000000"; 
      when 5325 => DO <= x"00000000"; 
      when 5326 => DO <= x"00000000"; 
      when 5327 => DO <= x"00000000"; 
      when 5328 => DO <= x"00000000"; 
      when 5329 => DO <= x"00000000"; 
      when 5330 => DO <= x"00000000"; 
      when 5331 => DO <= x"00000000"; 
      when 5332 => DO <= x"00000000"; 
      when 5333 => DO <= x"00000000"; 
      when 5334 => DO <= x"00000000"; 
      when 5335 => DO <= x"00000000"; 
      when 5336 => DO <= x"00000000"; 
      when 5337 => DO <= x"00000000"; 
      when 5338 => DO <= x"00000000"; 
      when 5339 => DO <= x"00000000"; 
      when 5340 => DO <= x"00000000"; 
      when 5341 => DO <= x"00000000"; 
      when 5342 => DO <= x"00000000"; 
      when 5343 => DO <= x"00000000"; 
      when 5344 => DO <= x"00000000"; 
      when 5345 => DO <= x"00000000"; 
      when 5346 => DO <= x"00000000"; 
      when 5347 => DO <= x"00000000"; 
      when 5348 => DO <= x"00000000"; 
      when 5349 => DO <= x"00000000"; 
      when 5350 => DO <= x"00000000"; 
      when 5351 => DO <= x"00000000"; 
      when 5352 => DO <= x"00000000"; 
      when 5353 => DO <= x"00000000"; 
      when 5354 => DO <= x"00000000"; 
      when 5355 => DO <= x"00000000"; 
      when 5356 => DO <= x"00000000"; 
      when 5357 => DO <= x"00000000"; 
      when 5358 => DO <= x"00000000"; 
      when 5359 => DO <= x"00000000"; 
      when 5360 => DO <= x"00000000"; 
      when 5361 => DO <= x"00000000"; 
      when 5362 => DO <= x"00000000"; 
      when 5363 => DO <= x"00000000"; 
      when 5364 => DO <= x"00000000"; 
      when 5365 => DO <= x"00000000"; 
      when 5366 => DO <= x"00000000"; 
      when 5367 => DO <= x"00000000"; 
      when 5368 => DO <= x"00000000"; 
      when 5369 => DO <= x"00000000"; 
      when 5370 => DO <= x"00000000"; 
      when 5371 => DO <= x"00000000"; 
      when 5372 => DO <= x"00000000"; 
      when 5373 => DO <= x"00000000"; 
      when 5374 => DO <= x"00000000"; 
      when 5375 => DO <= x"00000000"; 
      when 5376 => DO <= x"00000000"; 
      when 5377 => DO <= x"00000000"; 
      when 5378 => DO <= x"00000000"; 
      when 5379 => DO <= x"00000000"; 
      when 5380 => DO <= x"00000000"; 
      when 5381 => DO <= x"00000000"; 
      when 5382 => DO <= x"00000000"; 
      when 5383 => DO <= x"00000000"; 
      when 5384 => DO <= x"00000000"; 
      when 5385 => DO <= x"00000000"; 
      when 5386 => DO <= x"00000000"; 
      when 5387 => DO <= x"00000000"; 
      when 5388 => DO <= x"00000000"; 
      when 5389 => DO <= x"00000000"; 
      when 5390 => DO <= x"00000000"; 
      when 5391 => DO <= x"00000000"; 
      when 5392 => DO <= x"00000000"; 
      when 5393 => DO <= x"00000000"; 
      when 5394 => DO <= x"00000000"; 
      when 5395 => DO <= x"00000000"; 
      when 5396 => DO <= x"00000000"; 
      when 5397 => DO <= x"00000000"; 
      when 5398 => DO <= x"00000000"; 
      when 5399 => DO <= x"00000000"; 
      when 5400 => DO <= x"00000000"; 
      when 5401 => DO <= x"00000000"; 
      when 5402 => DO <= x"00000000"; 
      when 5403 => DO <= x"00000000"; 
      when 5404 => DO <= x"00000000"; 
      when 5405 => DO <= x"00000000"; 
      when 5406 => DO <= x"00000000"; 
      when 5407 => DO <= x"00000000"; 
      when 5408 => DO <= x"00000000"; 
      when 5409 => DO <= x"00000000"; 
      when 5410 => DO <= x"00000000"; 
      when 5411 => DO <= x"00000000"; 
      when 5412 => DO <= x"00000000"; 
      when 5413 => DO <= x"00000000"; 
      when 5414 => DO <= x"00000000"; 
      when 5415 => DO <= x"00000000"; 
      when 5416 => DO <= x"00000000"; 
      when 5417 => DO <= x"00000000"; 
      when 5418 => DO <= x"00000000"; 
      when 5419 => DO <= x"00000000"; 
      when 5420 => DO <= x"00000000"; 
      when 5421 => DO <= x"00000000"; 
      when 5422 => DO <= x"00000000"; 
      when 5423 => DO <= x"00000000"; 
      when 5424 => DO <= x"00000000"; 
      when 5425 => DO <= x"00000000"; 
      when 5426 => DO <= x"00000000"; 
      when 5427 => DO <= x"00000000"; 
      when 5428 => DO <= x"00000000"; 
      when 5429 => DO <= x"00000000"; 
      when 5430 => DO <= x"00000000"; 
      when 5431 => DO <= x"00000000"; 
      when 5432 => DO <= x"00000000"; 
      when 5433 => DO <= x"00000000"; 
      when 5434 => DO <= x"00000000"; 
      when 5435 => DO <= x"00000000"; 
      when 5436 => DO <= x"00000000"; 
      when 5437 => DO <= x"00000000"; 
      when 5438 => DO <= x"00000000"; 
      when 5439 => DO <= x"00000000"; 
      when 5440 => DO <= x"00000000"; 
      when 5441 => DO <= x"00000000"; 
      when 5442 => DO <= x"00000000"; 
      when 5443 => DO <= x"00000000"; 
      when 5444 => DO <= x"00000000"; 
      when 5445 => DO <= x"00000000"; 
      when 5446 => DO <= x"00000000"; 
      when 5447 => DO <= x"00000000"; 
      when 5448 => DO <= x"00000000"; 
      when 5449 => DO <= x"00000000"; 
      when 5450 => DO <= x"00000000"; 
      when 5451 => DO <= x"00000000"; 
      when 5452 => DO <= x"00000000"; 
      when 5453 => DO <= x"00000000"; 
      when 5454 => DO <= x"00000000"; 
      when 5455 => DO <= x"00000000"; 
      when 5456 => DO <= x"00000000"; 
      when 5457 => DO <= x"00000000"; 
      when 5458 => DO <= x"00000000"; 
      when 5459 => DO <= x"00000000"; 
      when 5460 => DO <= x"00000000"; 
      when 5461 => DO <= x"00000000"; 
      when 5462 => DO <= x"00000000"; 
      when 5463 => DO <= x"00000000"; 
      when 5464 => DO <= x"00000000"; 
      when 5465 => DO <= x"00000000"; 
      when 5466 => DO <= x"00000000"; 
      when 5467 => DO <= x"00000000"; 
      when 5468 => DO <= x"00000000"; 
      when 5469 => DO <= x"00000000"; 
      when 5470 => DO <= x"00000000"; 
      when 5471 => DO <= x"00000000"; 
      when 5472 => DO <= x"00000000"; 
      when 5473 => DO <= x"00000000"; 
      when 5474 => DO <= x"00000000"; 
      when 5475 => DO <= x"00000000"; 
      when 5476 => DO <= x"00000000"; 
      when 5477 => DO <= x"00000000"; 
      when 5478 => DO <= x"00000000"; 
      when 5479 => DO <= x"00000000"; 
      when 5480 => DO <= x"00000000"; 
      when 5481 => DO <= x"00000000"; 
      when 5482 => DO <= x"00000000"; 
      when 5483 => DO <= x"00000000"; 
      when 5484 => DO <= x"00000000"; 
      when 5485 => DO <= x"00000000"; 
      when 5486 => DO <= x"00000000"; 
      when 5487 => DO <= x"00000000"; 
      when 5488 => DO <= x"00000000"; 
      when 5489 => DO <= x"00000000"; 
      when 5490 => DO <= x"00000000"; 
      when 5491 => DO <= x"00000000"; 
      when 5492 => DO <= x"00000000"; 
      when 5493 => DO <= x"00000000"; 
      when 5494 => DO <= x"00000000"; 
      when 5495 => DO <= x"00000000"; 
      when 5496 => DO <= x"00000000"; 
      when 5497 => DO <= x"00000000"; 
      when 5498 => DO <= x"00000000"; 
      when 5499 => DO <= x"00000000"; 
      when 5500 => DO <= x"00000000"; 
      when 5501 => DO <= x"00000000"; 
      when 5502 => DO <= x"00000000"; 
      when 5503 => DO <= x"00000000"; 
      when 5504 => DO <= x"00000000"; 
      when 5505 => DO <= x"00000000"; 
      when 5506 => DO <= x"00000000"; 
      when 5507 => DO <= x"00000000"; 
      when 5508 => DO <= x"00000000"; 
      when 5509 => DO <= x"00000000"; 
      when 5510 => DO <= x"00000000"; 
      when 5511 => DO <= x"00000000"; 
      when 5512 => DO <= x"00000000"; 
      when 5513 => DO <= x"00000000"; 
      when 5514 => DO <= x"00000000"; 
      when 5515 => DO <= x"00000000"; 
      when 5516 => DO <= x"00000000"; 
      when 5517 => DO <= x"00000000"; 
      when 5518 => DO <= x"00000000"; 
      when 5519 => DO <= x"00000000"; 
      when 5520 => DO <= x"00000000"; 
      when 5521 => DO <= x"00000000"; 
      when 5522 => DO <= x"00000000"; 
      when 5523 => DO <= x"00000000"; 
      when 5524 => DO <= x"00000000"; 
      when 5525 => DO <= x"00000000"; 
      when 5526 => DO <= x"00000000"; 
      when 5527 => DO <= x"00000000"; 
      when 5528 => DO <= x"00000000"; 
      when 5529 => DO <= x"00000000"; 
      when 5530 => DO <= x"00000000"; 
      when 5531 => DO <= x"00000000"; 
      when 5532 => DO <= x"00000000"; 
      when 5533 => DO <= x"00000000"; 
      when 5534 => DO <= x"00000000"; 
      when 5535 => DO <= x"00000000"; 
      when 5536 => DO <= x"00000000"; 
      when 5537 => DO <= x"00000000"; 
      when 5538 => DO <= x"00000000"; 
      when 5539 => DO <= x"00000000"; 
      when 5540 => DO <= x"00000000"; 
      when 5541 => DO <= x"00000000"; 
      when 5542 => DO <= x"00000000"; 
      when 5543 => DO <= x"00000000"; 
      when 5544 => DO <= x"00000000"; 
      when 5545 => DO <= x"00000000"; 
      when 5546 => DO <= x"00000000"; 
      when 5547 => DO <= x"00000000"; 
      when 5548 => DO <= x"00000000"; 
      when 5549 => DO <= x"00000000"; 
      when 5550 => DO <= x"00000000"; 
      when 5551 => DO <= x"00000000"; 
      when 5552 => DO <= x"00000000"; 
      when 5553 => DO <= x"00000000"; 
      when 5554 => DO <= x"00000000"; 
      when 5555 => DO <= x"00000000"; 
      when 5556 => DO <= x"00000000"; 
      when 5557 => DO <= x"00000000"; 
      when 5558 => DO <= x"00000000"; 
      when 5559 => DO <= x"00000000"; 
      when 5560 => DO <= x"00000000"; 
      when 5561 => DO <= x"00000000"; 
      when 5562 => DO <= x"00000000"; 
      when 5563 => DO <= x"00000000"; 
      when 5564 => DO <= x"00000000"; 
      when 5565 => DO <= x"00000000"; 
      when 5566 => DO <= x"00000000"; 
      when 5567 => DO <= x"00000000"; 
      when 5568 => DO <= x"00000000"; 
      when 5569 => DO <= x"00000000"; 
      when 5570 => DO <= x"00000000"; 
      when 5571 => DO <= x"00000000"; 
      when 5572 => DO <= x"00000000"; 
      when 5573 => DO <= x"00000000"; 
      when 5574 => DO <= x"00000000"; 
      when 5575 => DO <= x"00000000"; 
      when 5576 => DO <= x"00000000"; 
      when 5577 => DO <= x"00000000"; 
      when 5578 => DO <= x"00000000"; 
      when 5579 => DO <= x"00000000"; 
      when 5580 => DO <= x"00000000"; 
      when 5581 => DO <= x"00000000"; 
      when 5582 => DO <= x"00000000"; 
      when 5583 => DO <= x"00000000"; 
      when 5584 => DO <= x"00000000"; 
      when 5585 => DO <= x"00000000"; 
      when 5586 => DO <= x"00000000"; 
      when 5587 => DO <= x"00000000"; 
      when 5588 => DO <= x"00000000"; 
      when 5589 => DO <= x"00000000"; 
      when 5590 => DO <= x"00000000"; 
      when 5591 => DO <= x"00000000"; 
      when 5592 => DO <= x"00000000"; 
      when 5593 => DO <= x"00000000"; 
      when 5594 => DO <= x"00000000"; 
      when 5595 => DO <= x"00000000"; 
      when 5596 => DO <= x"00000000"; 
      when 5597 => DO <= x"00000000"; 
      when 5598 => DO <= x"00000000"; 
      when 5599 => DO <= x"00000000"; 
      when 5600 => DO <= x"00000000"; 
      when 5601 => DO <= x"00000000"; 
      when 5602 => DO <= x"00000000"; 
      when 5603 => DO <= x"00000000"; 
      when 5604 => DO <= x"00000000"; 
      when 5605 => DO <= x"00000000"; 
      when 5606 => DO <= x"00000000"; 
      when 5607 => DO <= x"00000000"; 
      when 5608 => DO <= x"00000000"; 
      when 5609 => DO <= x"00000000"; 
      when 5610 => DO <= x"00000000"; 
      when 5611 => DO <= x"00000000"; 
      when 5612 => DO <= x"00000000"; 
      when 5613 => DO <= x"00000000"; 
      when 5614 => DO <= x"00000000"; 
      when 5615 => DO <= x"00000000"; 
      when 5616 => DO <= x"00000000"; 
      when 5617 => DO <= x"00000000"; 
      when 5618 => DO <= x"00000000"; 
      when 5619 => DO <= x"00000000"; 
      when 5620 => DO <= x"00000000"; 
      when 5621 => DO <= x"00000000"; 
      when 5622 => DO <= x"00000000"; 
      when 5623 => DO <= x"00000000"; 
      when 5624 => DO <= x"00000000"; 
      when 5625 => DO <= x"00000000"; 
      when 5626 => DO <= x"00000000"; 
      when 5627 => DO <= x"00000000"; 
      when 5628 => DO <= x"00000000"; 
      when 5629 => DO <= x"00000000"; 
      when 5630 => DO <= x"00000000"; 
      when 5631 => DO <= x"00000000"; 
      when 5632 => DO <= x"00000000"; 
      when 5633 => DO <= x"00000000"; 
      when 5634 => DO <= x"00000000"; 
      when 5635 => DO <= x"00000000"; 
      when 5636 => DO <= x"00000000"; 
      when 5637 => DO <= x"00000000"; 
      when 5638 => DO <= x"00000000"; 
      when 5639 => DO <= x"00000000"; 
      when 5640 => DO <= x"00000000"; 
      when 5641 => DO <= x"00000000"; 
      when 5642 => DO <= x"00000000"; 
      when 5643 => DO <= x"00000000"; 
      when 5644 => DO <= x"00000000"; 
      when 5645 => DO <= x"00000000"; 
      when 5646 => DO <= x"00000000"; 
      when 5647 => DO <= x"00000000"; 
      when 5648 => DO <= x"00000000"; 
      when 5649 => DO <= x"00000000"; 
      when 5650 => DO <= x"00000000"; 
      when 5651 => DO <= x"00000000"; 
      when 5652 => DO <= x"00000000"; 
      when 5653 => DO <= x"00000000"; 
      when 5654 => DO <= x"00000000"; 
      when 5655 => DO <= x"00000000"; 
      when 5656 => DO <= x"00000000"; 
      when 5657 => DO <= x"00000000"; 
      when 5658 => DO <= x"00000000"; 
      when 5659 => DO <= x"00000000"; 
      when 5660 => DO <= x"00000000"; 
      when 5661 => DO <= x"00000000"; 
      when 5662 => DO <= x"00000000"; 
      when 5663 => DO <= x"00000000"; 
      when 5664 => DO <= x"00000000"; 
      when 5665 => DO <= x"00000000"; 
      when 5666 => DO <= x"00000000"; 
      when 5667 => DO <= x"00000000"; 
      when 5668 => DO <= x"00000000"; 
      when 5669 => DO <= x"00000000"; 
      when 5670 => DO <= x"00000000"; 
      when 5671 => DO <= x"00000000"; 
      when 5672 => DO <= x"00000000"; 
      when 5673 => DO <= x"00000000"; 
      when 5674 => DO <= x"00000000"; 
      when 5675 => DO <= x"00000000"; 
      when 5676 => DO <= x"00000000"; 
      when 5677 => DO <= x"00000000"; 
      when 5678 => DO <= x"00000000"; 
      when 5679 => DO <= x"00000000"; 
      when 5680 => DO <= x"00000000"; 
      when 5681 => DO <= x"00000000"; 
      when 5682 => DO <= x"00000000"; 
      when 5683 => DO <= x"00000000"; 
      when 5684 => DO <= x"00000000"; 
      when 5685 => DO <= x"00000000"; 
      when 5686 => DO <= x"00000000"; 
      when 5687 => DO <= x"00000000"; 
      when 5688 => DO <= x"00000000"; 
      when 5689 => DO <= x"00000000"; 
      when 5690 => DO <= x"00000000"; 
      when 5691 => DO <= x"00000000"; 
      when 5692 => DO <= x"00000000"; 
      when 5693 => DO <= x"00000000"; 
      when 5694 => DO <= x"00000000"; 
      when 5695 => DO <= x"00000000"; 
      when 5696 => DO <= x"00000000"; 
      when 5697 => DO <= x"00000000"; 
      when 5698 => DO <= x"00000000"; 
      when 5699 => DO <= x"00000000"; 
      when 5700 => DO <= x"00000000"; 
      when 5701 => DO <= x"00000000"; 
      when 5702 => DO <= x"00000000"; 
      when 5703 => DO <= x"00000000"; 
      when 5704 => DO <= x"00000000"; 
      when 5705 => DO <= x"00000000"; 
      when 5706 => DO <= x"00000000"; 
      when 5707 => DO <= x"00000000"; 
      when 5708 => DO <= x"00000000"; 
      when 5709 => DO <= x"00000000"; 
      when 5710 => DO <= x"00000000"; 
      when 5711 => DO <= x"00000000"; 
      when 5712 => DO <= x"00000000"; 
      when 5713 => DO <= x"00000000"; 
      when 5714 => DO <= x"00000000"; 
      when 5715 => DO <= x"00000000"; 
      when 5716 => DO <= x"00000000"; 
      when 5717 => DO <= x"00000000"; 
      when 5718 => DO <= x"00000000"; 
      when 5719 => DO <= x"00000000"; 
      when 5720 => DO <= x"00000000"; 
      when 5721 => DO <= x"00000000"; 
      when 5722 => DO <= x"00000000"; 
      when 5723 => DO <= x"00000000"; 
      when 5724 => DO <= x"00000000"; 
      when 5725 => DO <= x"00000000"; 
      when 5726 => DO <= x"00000000"; 
      when 5727 => DO <= x"00000000"; 
      when 5728 => DO <= x"00000000"; 
      when 5729 => DO <= x"00000000"; 
      when 5730 => DO <= x"00000000"; 
      when 5731 => DO <= x"00000000"; 
      when 5732 => DO <= x"00000000"; 
      when 5733 => DO <= x"00000000"; 
      when 5734 => DO <= x"00000000"; 
      when 5735 => DO <= x"00000000"; 
      when 5736 => DO <= x"00000000"; 
      when 5737 => DO <= x"00000000"; 
      when 5738 => DO <= x"00000000"; 
      when 5739 => DO <= x"00000000"; 
      when 5740 => DO <= x"00000000"; 
      when 5741 => DO <= x"00000000"; 
      when 5742 => DO <= x"00000000"; 
      when 5743 => DO <= x"00000000"; 
      when 5744 => DO <= x"00000000"; 
      when 5745 => DO <= x"00000000"; 
      when 5746 => DO <= x"00000000"; 
      when 5747 => DO <= x"00000000"; 
      when 5748 => DO <= x"00000000"; 
      when 5749 => DO <= x"00000000"; 
      when 5750 => DO <= x"00000000"; 
      when 5751 => DO <= x"00000000"; 
      when 5752 => DO <= x"00000000"; 
      when 5753 => DO <= x"00000000"; 
      when 5754 => DO <= x"00000000"; 
      when 5755 => DO <= x"00000000"; 
      when 5756 => DO <= x"00000000"; 
      when 5757 => DO <= x"00000000"; 
      when 5758 => DO <= x"00000000"; 
      when 5759 => DO <= x"00000000"; 
      when 5760 => DO <= x"00000000"; 
      when 5761 => DO <= x"00000000"; 
      when 5762 => DO <= x"00000000"; 
      when 5763 => DO <= x"00000000"; 
      when 5764 => DO <= x"00000000"; 
      when 5765 => DO <= x"00000000"; 
      when 5766 => DO <= x"00000000"; 
      when 5767 => DO <= x"00000000"; 
      when 5768 => DO <= x"00000000"; 
      when 5769 => DO <= x"00000000"; 
      when 5770 => DO <= x"00000000"; 
      when 5771 => DO <= x"00000000"; 
      when 5772 => DO <= x"00000000"; 
      when 5773 => DO <= x"00000000"; 
      when 5774 => DO <= x"00000000"; 
      when 5775 => DO <= x"00000000"; 
      when 5776 => DO <= x"00000000"; 
      when 5777 => DO <= x"00000000"; 
      when 5778 => DO <= x"00000000"; 
      when 5779 => DO <= x"00000000"; 
      when 5780 => DO <= x"00000000"; 
      when 5781 => DO <= x"00000000"; 
      when 5782 => DO <= x"00000000"; 
      when 5783 => DO <= x"00000000"; 
      when 5784 => DO <= x"00000000"; 
      when 5785 => DO <= x"00000000"; 
      when 5786 => DO <= x"00000000"; 
      when 5787 => DO <= x"00000000"; 
      when 5788 => DO <= x"00000000"; 
      when 5789 => DO <= x"00000000"; 
      when 5790 => DO <= x"00000000"; 
      when 5791 => DO <= x"00000000"; 
      when 5792 => DO <= x"00000000"; 
      when 5793 => DO <= x"00000000"; 
      when 5794 => DO <= x"00000000"; 
      when 5795 => DO <= x"00000000"; 
      when 5796 => DO <= x"00000000"; 
      when 5797 => DO <= x"00000000"; 
      when 5798 => DO <= x"00000000"; 
      when 5799 => DO <= x"00000000"; 
      when 5800 => DO <= x"00000000"; 
      when 5801 => DO <= x"00000000"; 
      when 5802 => DO <= x"00000000"; 
      when 5803 => DO <= x"00000000"; 
      when 5804 => DO <= x"00000000"; 
      when 5805 => DO <= x"00000000"; 
      when 5806 => DO <= x"00000000"; 
      when 5807 => DO <= x"00000000"; 
      when 5808 => DO <= x"00000000"; 
      when 5809 => DO <= x"00000000"; 
      when 5810 => DO <= x"00000000"; 
      when 5811 => DO <= x"00000000"; 
      when 5812 => DO <= x"00000000"; 
      when 5813 => DO <= x"00000000"; 
      when 5814 => DO <= x"00000000"; 
      when 5815 => DO <= x"00000000"; 
      when 5816 => DO <= x"00000000"; 
      when 5817 => DO <= x"00000000"; 
      when 5818 => DO <= x"00000000"; 
      when 5819 => DO <= x"00000000"; 
      when 5820 => DO <= x"00000000"; 
      when 5821 => DO <= x"00000000"; 
      when 5822 => DO <= x"00000000"; 
      when 5823 => DO <= x"00000000"; 
      when 5824 => DO <= x"00000000"; 
      when 5825 => DO <= x"00000000"; 
      when 5826 => DO <= x"00000000"; 
      when 5827 => DO <= x"00000000"; 
      when 5828 => DO <= x"00000000"; 
      when 5829 => DO <= x"00000000"; 
      when 5830 => DO <= x"00000000"; 
      when 5831 => DO <= x"00000000"; 
      when 5832 => DO <= x"00000000"; 
      when 5833 => DO <= x"00000000"; 
      when 5834 => DO <= x"00000000"; 
      when 5835 => DO <= x"00000000"; 
      when 5836 => DO <= x"00000000"; 
      when 5837 => DO <= x"00000000"; 
      when 5838 => DO <= x"00000000"; 
      when 5839 => DO <= x"00000000"; 
      when 5840 => DO <= x"00000000"; 
      when 5841 => DO <= x"00000000"; 
      when 5842 => DO <= x"00000000"; 
      when 5843 => DO <= x"00000000"; 
      when 5844 => DO <= x"00000000"; 
      when 5845 => DO <= x"00000000"; 
      when 5846 => DO <= x"00000000"; 
      when 5847 => DO <= x"00000000"; 
      when 5848 => DO <= x"00000000"; 
      when 5849 => DO <= x"00000000"; 
      when 5850 => DO <= x"00000000"; 
      when 5851 => DO <= x"00000000"; 
      when 5852 => DO <= x"00000000"; 
      when 5853 => DO <= x"00000000"; 
      when 5854 => DO <= x"00000000"; 
      when 5855 => DO <= x"00000000"; 
      when 5856 => DO <= x"00000000"; 
      when 5857 => DO <= x"00000000"; 
      when 5858 => DO <= x"00000000"; 
      when 5859 => DO <= x"00000000"; 
      when 5860 => DO <= x"00000000"; 
      when 5861 => DO <= x"00000000"; 
      when 5862 => DO <= x"00000000"; 
      when 5863 => DO <= x"00000000"; 
      when 5864 => DO <= x"00000000"; 
      when 5865 => DO <= x"00000000"; 
      when 5866 => DO <= x"00000000"; 
      when 5867 => DO <= x"00000000"; 
      when 5868 => DO <= x"00000000"; 
      when 5869 => DO <= x"00000000"; 
      when 5870 => DO <= x"00000000"; 
      when 5871 => DO <= x"00000000"; 
      when 5872 => DO <= x"00000000"; 
      when 5873 => DO <= x"00000000"; 
      when 5874 => DO <= x"00000000"; 
      when 5875 => DO <= x"00000000"; 
      when 5876 => DO <= x"00000000"; 
      when 5877 => DO <= x"00000000"; 
      when 5878 => DO <= x"00000000"; 
      when 5879 => DO <= x"00000000"; 
      when 5880 => DO <= x"00000000"; 
      when 5881 => DO <= x"00000000"; 
      when 5882 => DO <= x"00000000"; 
      when 5883 => DO <= x"00000000"; 
      when 5884 => DO <= x"00000000"; 
      when 5885 => DO <= x"00000000"; 
      when 5886 => DO <= x"00000000"; 
      when 5887 => DO <= x"00000000"; 
      when 5888 => DO <= x"00000000"; 
      when 5889 => DO <= x"00000000"; 
      when 5890 => DO <= x"00000000"; 
      when 5891 => DO <= x"00000000"; 
      when 5892 => DO <= x"00000000"; 
      when 5893 => DO <= x"00000000"; 
      when 5894 => DO <= x"00000000"; 
      when 5895 => DO <= x"00000000"; 
      when 5896 => DO <= x"00000000"; 
      when 5897 => DO <= x"00000000"; 
      when 5898 => DO <= x"00000000"; 
      when 5899 => DO <= x"00000000"; 
      when 5900 => DO <= x"00000000"; 
      when 5901 => DO <= x"00000000"; 
      when 5902 => DO <= x"00000000"; 
      when 5903 => DO <= x"00000000"; 
      when 5904 => DO <= x"00000000"; 
      when 5905 => DO <= x"00000000"; 
      when 5906 => DO <= x"00000000"; 
      when 5907 => DO <= x"00000000"; 
      when 5908 => DO <= x"00000000"; 
      when 5909 => DO <= x"00000000"; 
      when 5910 => DO <= x"00000000"; 
      when 5911 => DO <= x"00000000"; 
      when 5912 => DO <= x"00000000"; 
      when 5913 => DO <= x"00000000"; 
      when 5914 => DO <= x"00000000"; 
      when 5915 => DO <= x"00000000"; 
      when 5916 => DO <= x"00000000"; 
      when 5917 => DO <= x"00000000"; 
      when 5918 => DO <= x"00000000"; 
      when 5919 => DO <= x"00000000"; 
      when 5920 => DO <= x"00000000"; 
      when 5921 => DO <= x"00000000"; 
      when 5922 => DO <= x"00000000"; 
      when 5923 => DO <= x"00000000"; 
      when 5924 => DO <= x"00000000"; 
      when 5925 => DO <= x"00000000"; 
      when 5926 => DO <= x"00000000"; 
      when 5927 => DO <= x"00000000"; 
      when 5928 => DO <= x"00000000"; 
      when 5929 => DO <= x"00000000"; 
      when 5930 => DO <= x"00000000"; 
      when 5931 => DO <= x"00000000"; 
      when 5932 => DO <= x"00000000"; 
      when 5933 => DO <= x"00000000"; 
      when 5934 => DO <= x"00000000"; 
      when 5935 => DO <= x"00000000"; 
      when 5936 => DO <= x"00000000"; 
      when 5937 => DO <= x"00000000"; 
      when 5938 => DO <= x"00000000"; 
      when 5939 => DO <= x"00000000"; 
      when 5940 => DO <= x"00000000"; 
      when 5941 => DO <= x"00000000"; 
      when 5942 => DO <= x"00000000"; 
      when 5943 => DO <= x"00000000"; 
      when 5944 => DO <= x"00000000"; 
      when 5945 => DO <= x"00000000"; 
      when 5946 => DO <= x"00000000"; 
      when 5947 => DO <= x"00000000"; 
      when 5948 => DO <= x"00000000"; 
      when 5949 => DO <= x"00000000"; 
      when 5950 => DO <= x"00000000"; 
      when 5951 => DO <= x"00000000"; 
      when 5952 => DO <= x"00000000"; 
      when 5953 => DO <= x"00000000"; 
      when 5954 => DO <= x"00000000"; 
      when 5955 => DO <= x"00000000"; 
      when 5956 => DO <= x"00000000"; 
      when 5957 => DO <= x"00000000"; 
      when 5958 => DO <= x"00000000"; 
      when 5959 => DO <= x"00000000"; 
      when 5960 => DO <= x"00000000"; 
      when 5961 => DO <= x"00000000"; 
      when 5962 => DO <= x"00000000"; 
      when 5963 => DO <= x"00000000"; 
      when 5964 => DO <= x"00000000"; 
      when 5965 => DO <= x"00000000"; 
      when 5966 => DO <= x"00000000"; 
      when 5967 => DO <= x"00000000"; 
      when 5968 => DO <= x"00000000"; 
      when 5969 => DO <= x"00000000"; 
      when 5970 => DO <= x"00000000"; 
      when 5971 => DO <= x"00000000"; 
      when 5972 => DO <= x"00000000"; 
      when 5973 => DO <= x"00000000"; 
      when 5974 => DO <= x"00000000"; 
      when 5975 => DO <= x"00000000"; 
      when 5976 => DO <= x"00000000"; 
      when 5977 => DO <= x"00000000"; 
      when 5978 => DO <= x"00000000"; 
      when 5979 => DO <= x"00000000"; 
      when 5980 => DO <= x"00000000"; 
      when 5981 => DO <= x"00000000"; 
      when 5982 => DO <= x"00000000"; 
      when 5983 => DO <= x"00000000"; 
      when 5984 => DO <= x"00000000"; 
      when 5985 => DO <= x"00000000"; 
      when 5986 => DO <= x"00000000"; 
      when 5987 => DO <= x"00000000"; 
      when 5988 => DO <= x"00000000"; 
      when 5989 => DO <= x"00000000"; 
      when 5990 => DO <= x"00000000"; 
      when 5991 => DO <= x"00000000"; 
      when 5992 => DO <= x"00000000"; 
      when 5993 => DO <= x"00000000"; 
      when 5994 => DO <= x"00000000"; 
      when 5995 => DO <= x"00000000"; 
      when 5996 => DO <= x"00000000"; 
      when 5997 => DO <= x"00000000"; 
      when 5998 => DO <= x"00000000"; 
      when 5999 => DO <= x"00000000"; 
      when 6000 => DO <= x"00000000"; 
      when 6001 => DO <= x"00000000"; 
      when 6002 => DO <= x"00000000"; 
      when 6003 => DO <= x"00000000"; 
      when 6004 => DO <= x"00000000"; 
      when 6005 => DO <= x"00000000"; 
      when 6006 => DO <= x"00000000"; 
      when 6007 => DO <= x"00000000"; 
      when 6008 => DO <= x"00000000"; 
      when 6009 => DO <= x"00000000"; 
      when 6010 => DO <= x"00000000"; 
      when 6011 => DO <= x"00000000"; 
      when 6012 => DO <= x"00000000"; 
      when 6013 => DO <= x"00000000"; 
      when 6014 => DO <= x"00000000"; 
      when 6015 => DO <= x"00000000"; 
      when 6016 => DO <= x"00000000"; 
      when 6017 => DO <= x"00000000"; 
      when 6018 => DO <= x"00000000"; 
      when 6019 => DO <= x"00000000"; 
      when 6020 => DO <= x"00000000"; 
      when 6021 => DO <= x"00000000"; 
      when 6022 => DO <= x"00000000"; 
      when 6023 => DO <= x"00000000"; 
      when 6024 => DO <= x"00000000"; 
      when 6025 => DO <= x"00000000"; 
      when 6026 => DO <= x"00000000"; 
      when 6027 => DO <= x"00000000"; 
      when 6028 => DO <= x"00000000"; 
      when 6029 => DO <= x"00000000"; 
      when 6030 => DO <= x"00000000"; 
      when 6031 => DO <= x"00000000"; 
      when 6032 => DO <= x"00000000"; 
      when 6033 => DO <= x"00000000"; 
      when 6034 => DO <= x"00000000"; 
      when 6035 => DO <= x"00000000"; 
      when 6036 => DO <= x"00000000"; 
      when 6037 => DO <= x"00000000"; 
      when 6038 => DO <= x"00000000"; 
      when 6039 => DO <= x"00000000"; 
      when 6040 => DO <= x"00000000"; 
      when 6041 => DO <= x"00000000"; 
      when 6042 => DO <= x"00000000"; 
      when 6043 => DO <= x"00000000"; 
      when 6044 => DO <= x"00000000"; 
      when 6045 => DO <= x"00000000"; 
      when 6046 => DO <= x"00000000"; 
      when 6047 => DO <= x"00000000"; 
      when 6048 => DO <= x"00000000"; 
      when 6049 => DO <= x"00000000"; 
      when 6050 => DO <= x"00000000"; 
      when 6051 => DO <= x"00000000"; 
      when 6052 => DO <= x"00000000"; 
      when 6053 => DO <= x"00000000"; 
      when 6054 => DO <= x"00000000"; 
      when 6055 => DO <= x"00000000"; 
      when 6056 => DO <= x"00000000"; 
      when 6057 => DO <= x"00000000"; 
      when 6058 => DO <= x"00000000"; 
      when 6059 => DO <= x"00000000"; 
      when 6060 => DO <= x"00000000"; 
      when 6061 => DO <= x"00000000"; 
      when 6062 => DO <= x"00000000"; 
      when 6063 => DO <= x"00000000"; 
      when 6064 => DO <= x"00000000"; 
      when 6065 => DO <= x"00000000"; 
      when 6066 => DO <= x"00000000"; 
      when 6067 => DO <= x"00000000"; 
      when 6068 => DO <= x"00000000"; 
      when 6069 => DO <= x"00000000"; 
      when 6070 => DO <= x"00000000"; 
      when 6071 => DO <= x"00000000"; 
      when 6072 => DO <= x"00000000"; 
      when 6073 => DO <= x"00000000"; 
      when 6074 => DO <= x"00000000"; 
      when 6075 => DO <= x"00000000"; 
      when 6076 => DO <= x"00000000"; 
      when 6077 => DO <= x"00000000"; 
      when 6078 => DO <= x"00000000"; 
      when 6079 => DO <= x"00000000"; 
      when 6080 => DO <= x"00000000"; 
      when 6081 => DO <= x"00000000"; 
      when 6082 => DO <= x"00000000"; 
      when 6083 => DO <= x"00000000"; 
      when 6084 => DO <= x"00000000"; 
      when 6085 => DO <= x"00000000"; 
      when 6086 => DO <= x"00000000"; 
      when 6087 => DO <= x"00000000"; 
      when 6088 => DO <= x"00000000"; 
      when 6089 => DO <= x"00000000"; 
      when 6090 => DO <= x"00000000"; 
      when 6091 => DO <= x"00000000"; 
      when 6092 => DO <= x"00000000"; 
      when 6093 => DO <= x"00000000"; 
      when 6094 => DO <= x"00000000"; 
      when 6095 => DO <= x"00000000"; 
      when 6096 => DO <= x"00000000"; 
      when 6097 => DO <= x"00000000"; 
      when 6098 => DO <= x"00000000"; 
      when 6099 => DO <= x"00000000"; 
      when 6100 => DO <= x"00000000"; 
      when 6101 => DO <= x"00000000"; 
      when 6102 => DO <= x"00000000"; 
      when 6103 => DO <= x"00000000"; 
      when 6104 => DO <= x"00000000"; 
      when 6105 => DO <= x"00000000"; 
      when 6106 => DO <= x"00000000"; 
      when 6107 => DO <= x"00000000"; 
      when 6108 => DO <= x"00000000"; 
      when 6109 => DO <= x"00000000"; 
      when 6110 => DO <= x"00000000"; 
      when 6111 => DO <= x"00000000"; 
      when 6112 => DO <= x"00000000"; 
      when 6113 => DO <= x"00000000"; 
      when 6114 => DO <= x"00000000"; 
      when 6115 => DO <= x"00000000"; 
      when 6116 => DO <= x"00000000"; 
      when 6117 => DO <= x"00000000"; 
      when 6118 => DO <= x"00000000"; 
      when 6119 => DO <= x"00000000"; 
      when 6120 => DO <= x"00000000"; 
      when 6121 => DO <= x"00000000"; 
      when 6122 => DO <= x"00000000"; 
      when 6123 => DO <= x"00000000"; 
      when 6124 => DO <= x"00000000"; 
      when 6125 => DO <= x"00000000"; 
      when 6126 => DO <= x"00000000"; 
      when 6127 => DO <= x"00000000"; 
      when 6128 => DO <= x"00000000"; 
      when 6129 => DO <= x"00000000"; 
      when 6130 => DO <= x"00000000"; 
      when 6131 => DO <= x"00000000"; 
      when 6132 => DO <= x"00000000"; 
      when 6133 => DO <= x"00000000"; 
      when 6134 => DO <= x"00000000"; 
      when 6135 => DO <= x"00000000"; 
      when 6136 => DO <= x"00000000"; 
      when 6137 => DO <= x"00000000"; 
      when 6138 => DO <= x"00000000"; 
      when 6139 => DO <= x"00000000"; 
      when 6140 => DO <= x"00000000"; 
      when 6141 => DO <= x"00000000"; 
      when 6142 => DO <= x"00000000"; 
      when 6143 => DO <= x"00000000"; 
      when 6144 => DO <= x"00000000"; 
      when 6145 => DO <= x"00000000"; 
      when 6146 => DO <= x"00000000"; 
      when 6147 => DO <= x"00000000"; 
      when 6148 => DO <= x"00000000"; 
      when 6149 => DO <= x"00000000"; 
      when 6150 => DO <= x"00000000"; 
      when 6151 => DO <= x"00000000"; 
      when 6152 => DO <= x"00000000"; 
      when 6153 => DO <= x"00000000"; 
      when 6154 => DO <= x"00000000"; 
      when 6155 => DO <= x"00000000"; 
      when 6156 => DO <= x"00000000"; 
      when 6157 => DO <= x"00000000"; 
      when 6158 => DO <= x"00000000"; 
      when 6159 => DO <= x"00000000"; 
      when 6160 => DO <= x"00000000"; 
      when 6161 => DO <= x"00000000"; 
      when 6162 => DO <= x"00000000"; 
      when 6163 => DO <= x"00000000"; 
      when 6164 => DO <= x"00000000"; 
      when 6165 => DO <= x"00000000"; 
      when 6166 => DO <= x"00000000"; 
      when 6167 => DO <= x"00000000"; 
      when 6168 => DO <= x"00000000"; 
      when 6169 => DO <= x"00000000"; 
      when 6170 => DO <= x"00000000"; 
      when 6171 => DO <= x"00000000"; 
      when 6172 => DO <= x"00000000"; 
      when 6173 => DO <= x"00000000"; 
      when 6174 => DO <= x"00000000"; 
      when 6175 => DO <= x"00000000"; 
      when 6176 => DO <= x"00000000"; 
      when 6177 => DO <= x"00000000"; 
      when 6178 => DO <= x"00000000"; 
      when 6179 => DO <= x"00000000"; 
      when 6180 => DO <= x"00000000"; 
      when 6181 => DO <= x"00000000"; 
      when 6182 => DO <= x"00000000"; 
      when 6183 => DO <= x"00000000"; 
      when 6184 => DO <= x"00000000"; 
      when 6185 => DO <= x"00000000"; 
      when 6186 => DO <= x"00000000"; 
      when 6187 => DO <= x"00000000"; 
      when 6188 => DO <= x"00000000"; 
      when 6189 => DO <= x"00000000"; 
      when 6190 => DO <= x"00000000"; 
      when 6191 => DO <= x"00000000"; 
      when 6192 => DO <= x"00000000"; 
      when 6193 => DO <= x"00000000"; 
      when 6194 => DO <= x"00000000"; 
      when 6195 => DO <= x"00000000"; 
      when 6196 => DO <= x"00000000"; 
      when 6197 => DO <= x"00000000"; 
      when 6198 => DO <= x"00000000"; 
      when 6199 => DO <= x"00000000"; 
      when 6200 => DO <= x"00000000"; 
      when 6201 => DO <= x"00000000"; 
      when 6202 => DO <= x"00000000"; 
      when 6203 => DO <= x"00000000"; 
      when 6204 => DO <= x"00000000"; 
      when 6205 => DO <= x"00000000"; 
      when 6206 => DO <= x"00000000"; 
      when 6207 => DO <= x"00000000"; 
      when 6208 => DO <= x"00000000"; 
      when 6209 => DO <= x"00000000"; 
      when 6210 => DO <= x"00000000"; 
      when 6211 => DO <= x"00000000"; 
      when 6212 => DO <= x"00000000"; 
      when 6213 => DO <= x"00000000"; 
      when 6214 => DO <= x"00000000"; 
      when 6215 => DO <= x"00000000"; 
      when 6216 => DO <= x"00000000"; 
      when 6217 => DO <= x"00000000"; 
      when 6218 => DO <= x"00000000"; 
      when 6219 => DO <= x"00000000"; 
      when 6220 => DO <= x"00000000"; 
      when 6221 => DO <= x"00000000"; 
      when 6222 => DO <= x"00000000"; 
      when 6223 => DO <= x"00000000"; 
      when 6224 => DO <= x"00000000"; 
      when 6225 => DO <= x"00000000"; 
      when 6226 => DO <= x"00000000"; 
      when 6227 => DO <= x"00000000"; 
      when 6228 => DO <= x"00000000"; 
      when 6229 => DO <= x"00000000"; 
      when 6230 => DO <= x"00000000"; 
      when 6231 => DO <= x"00000000"; 
      when 6232 => DO <= x"00000000"; 
      when 6233 => DO <= x"00000000"; 
      when 6234 => DO <= x"00000000"; 
      when 6235 => DO <= x"00000000"; 
      when 6236 => DO <= x"00000000"; 
      when 6237 => DO <= x"00000000"; 
      when 6238 => DO <= x"00000000"; 
      when 6239 => DO <= x"00000000"; 
      when 6240 => DO <= x"00000000"; 
      when 6241 => DO <= x"00000000"; 
      when 6242 => DO <= x"00000000"; 
      when 6243 => DO <= x"00000000"; 
      when 6244 => DO <= x"00000000"; 
      when 6245 => DO <= x"00000000"; 
      when 6246 => DO <= x"00000000"; 
      when 6247 => DO <= x"00000000"; 
      when 6248 => DO <= x"00000000"; 
      when 6249 => DO <= x"00000000"; 
      when 6250 => DO <= x"00000000"; 
      when 6251 => DO <= x"00000000"; 
      when 6252 => DO <= x"00000000"; 
      when 6253 => DO <= x"00000000"; 
      when 6254 => DO <= x"00000000"; 
      when 6255 => DO <= x"00000000"; 
      when 6256 => DO <= x"00000000"; 
      when 6257 => DO <= x"00000000"; 
      when 6258 => DO <= x"00000000"; 
      when 6259 => DO <= x"00000000"; 
      when 6260 => DO <= x"00000000"; 
      when 6261 => DO <= x"00000000"; 
      when 6262 => DO <= x"00000000"; 
      when 6263 => DO <= x"00000000"; 
      when 6264 => DO <= x"00000000"; 
      when 6265 => DO <= x"00000000"; 
      when 6266 => DO <= x"00000000"; 
      when 6267 => DO <= x"00000000"; 
      when 6268 => DO <= x"00000000"; 
      when 6269 => DO <= x"00000000"; 
      when 6270 => DO <= x"00000000"; 
      when 6271 => DO <= x"00000000"; 
      when 6272 => DO <= x"00000000"; 
      when 6273 => DO <= x"00000000"; 
      when 6274 => DO <= x"00000000"; 
      when 6275 => DO <= x"00000000"; 
      when 6276 => DO <= x"00000000"; 
      when 6277 => DO <= x"00000000"; 
      when 6278 => DO <= x"00000000"; 
      when 6279 => DO <= x"00000000"; 
      when 6280 => DO <= x"00000000"; 
      when 6281 => DO <= x"00000000"; 
      when 6282 => DO <= x"00000000"; 
      when 6283 => DO <= x"00000000"; 
      when 6284 => DO <= x"00000000"; 
      when 6285 => DO <= x"00000000"; 
      when 6286 => DO <= x"00000000"; 
      when 6287 => DO <= x"00000000"; 
      when 6288 => DO <= x"00000000"; 
      when 6289 => DO <= x"00000000"; 
      when 6290 => DO <= x"00000000"; 
      when 6291 => DO <= x"00000000"; 
      when 6292 => DO <= x"00000000"; 
      when 6293 => DO <= x"00000000"; 
      when 6294 => DO <= x"00000000"; 
      when 6295 => DO <= x"00000000"; 
      when 6296 => DO <= x"00000000"; 
      when 6297 => DO <= x"00000000"; 
      when 6298 => DO <= x"00000000"; 
      when 6299 => DO <= x"00000000"; 
      when 6300 => DO <= x"00000000"; 
      when 6301 => DO <= x"00000000"; 
      when 6302 => DO <= x"00000000"; 
      when 6303 => DO <= x"00000000"; 
      when 6304 => DO <= x"00000000"; 
      when 6305 => DO <= x"00000000"; 
      when 6306 => DO <= x"00000000"; 
      when 6307 => DO <= x"00000000"; 
      when 6308 => DO <= x"00000000"; 
      when 6309 => DO <= x"00000000"; 
      when 6310 => DO <= x"00000000"; 
      when 6311 => DO <= x"00000000"; 
      when 6312 => DO <= x"00000000"; 
      when 6313 => DO <= x"00000000"; 
      when 6314 => DO <= x"00000000"; 
      when 6315 => DO <= x"00000000"; 
      when 6316 => DO <= x"00000000"; 
      when 6317 => DO <= x"00000000"; 
      when 6318 => DO <= x"00000000"; 
      when 6319 => DO <= x"00000000"; 
      when 6320 => DO <= x"00000000"; 
      when 6321 => DO <= x"00000000"; 
      when 6322 => DO <= x"00000000"; 
      when 6323 => DO <= x"00000000"; 
      when 6324 => DO <= x"00000000"; 
      when 6325 => DO <= x"00000000"; 
      when 6326 => DO <= x"00000000"; 
      when 6327 => DO <= x"00000000"; 
      when 6328 => DO <= x"00000000"; 
      when 6329 => DO <= x"00000000"; 
      when 6330 => DO <= x"00000000"; 
      when 6331 => DO <= x"00000000"; 
      when 6332 => DO <= x"00000000"; 
      when 6333 => DO <= x"00000000"; 
      when 6334 => DO <= x"00000000"; 
      when 6335 => DO <= x"00000000"; 
      when 6336 => DO <= x"00000000"; 
      when 6337 => DO <= x"00000000"; 
      when 6338 => DO <= x"00000000"; 
      when 6339 => DO <= x"00000000"; 
      when 6340 => DO <= x"00000000"; 
      when 6341 => DO <= x"00000000"; 
      when 6342 => DO <= x"00000000"; 
      when 6343 => DO <= x"00000000"; 
      when 6344 => DO <= x"00000000"; 
      when 6345 => DO <= x"00000000"; 
      when 6346 => DO <= x"00000000"; 
      when 6347 => DO <= x"00000000"; 
      when 6348 => DO <= x"00000000"; 
      when 6349 => DO <= x"00000000"; 
      when 6350 => DO <= x"00000000"; 
      when 6351 => DO <= x"00000000"; 
      when 6352 => DO <= x"00000000"; 
      when 6353 => DO <= x"00000000"; 
      when 6354 => DO <= x"00000000"; 
      when 6355 => DO <= x"00000000"; 
      when 6356 => DO <= x"00000000"; 
      when 6357 => DO <= x"00000000"; 
      when 6358 => DO <= x"00000000"; 
      when 6359 => DO <= x"00000000"; 
      when 6360 => DO <= x"00000000"; 
      when 6361 => DO <= x"00000000"; 
      when 6362 => DO <= x"00000000"; 
      when 6363 => DO <= x"00000000"; 
      when 6364 => DO <= x"00000000"; 
      when 6365 => DO <= x"00000000"; 
      when 6366 => DO <= x"00000000"; 
      when 6367 => DO <= x"00000000"; 
      when 6368 => DO <= x"00000000"; 
      when 6369 => DO <= x"00000000"; 
      when 6370 => DO <= x"00000000"; 
      when 6371 => DO <= x"00000000"; 
      when 6372 => DO <= x"00000000"; 
      when 6373 => DO <= x"00000000"; 
      when 6374 => DO <= x"00000000"; 
      when 6375 => DO <= x"00000000"; 
      when 6376 => DO <= x"00000000"; 
      when 6377 => DO <= x"00000000"; 
      when 6378 => DO <= x"00000000"; 
      when 6379 => DO <= x"00000000"; 
      when 6380 => DO <= x"00000000"; 
      when 6381 => DO <= x"00000000"; 
      when 6382 => DO <= x"00000000"; 
      when 6383 => DO <= x"00000000"; 
      when 6384 => DO <= x"00000000"; 
      when 6385 => DO <= x"00000000"; 
      when 6386 => DO <= x"00000000"; 
      when 6387 => DO <= x"00000000"; 
      when 6388 => DO <= x"00000000"; 
      when 6389 => DO <= x"00000000"; 
      when 6390 => DO <= x"00000000"; 
      when 6391 => DO <= x"00000000"; 
      when 6392 => DO <= x"00000000"; 
      when 6393 => DO <= x"00000000"; 
      when 6394 => DO <= x"00000000"; 
      when 6395 => DO <= x"00000000"; 
      when 6396 => DO <= x"00000000"; 
      when 6397 => DO <= x"00000000"; 
      when 6398 => DO <= x"00000000"; 
      when 6399 => DO <= x"00000000"; 
      when 6400 => DO <= x"00000000"; 
      when 6401 => DO <= x"00000000"; 
      when 6402 => DO <= x"00000000"; 
      when 6403 => DO <= x"00000000"; 
      when 6404 => DO <= x"00000000"; 
      when 6405 => DO <= x"00000000"; 
      when 6406 => DO <= x"00000000"; 
      when 6407 => DO <= x"00000000"; 
      when 6408 => DO <= x"00000000"; 
      when 6409 => DO <= x"00000000"; 
      when 6410 => DO <= x"00000000"; 
      when 6411 => DO <= x"00000000"; 
      when 6412 => DO <= x"00000000"; 
      when 6413 => DO <= x"00000000"; 
      when 6414 => DO <= x"00000000"; 
      when 6415 => DO <= x"00000000"; 
      when 6416 => DO <= x"00000000"; 
      when 6417 => DO <= x"00000000"; 
      when 6418 => DO <= x"00000000"; 
      when 6419 => DO <= x"00000000"; 
      when 6420 => DO <= x"00000000"; 
      when 6421 => DO <= x"00000000"; 
      when 6422 => DO <= x"00000000"; 
      when 6423 => DO <= x"00000000"; 
      when 6424 => DO <= x"00000000"; 
      when 6425 => DO <= x"00000000"; 
      when 6426 => DO <= x"00000000"; 
      when 6427 => DO <= x"00000000"; 
      when 6428 => DO <= x"00000000"; 
      when 6429 => DO <= x"00000000"; 
      when 6430 => DO <= x"00000000"; 
      when 6431 => DO <= x"00000000"; 
      when 6432 => DO <= x"00000000"; 
      when 6433 => DO <= x"00000000"; 
      when 6434 => DO <= x"00000000"; 
      when 6435 => DO <= x"00000000"; 
      when 6436 => DO <= x"00000000"; 
      when 6437 => DO <= x"00000000"; 
      when 6438 => DO <= x"00000000"; 
      when 6439 => DO <= x"00000000"; 
      when 6440 => DO <= x"00000000"; 
      when 6441 => DO <= x"00000000"; 
      when 6442 => DO <= x"00000000"; 
      when 6443 => DO <= x"00000000"; 
      when 6444 => DO <= x"00000000"; 
      when 6445 => DO <= x"00000000"; 
      when 6446 => DO <= x"00000000"; 
      when 6447 => DO <= x"00000000"; 
      when 6448 => DO <= x"00000000"; 
      when 6449 => DO <= x"00000000"; 
      when 6450 => DO <= x"00000000"; 
      when 6451 => DO <= x"00000000"; 
      when 6452 => DO <= x"00000000"; 
      when 6453 => DO <= x"00000000"; 
      when 6454 => DO <= x"00000000"; 
      when 6455 => DO <= x"00000000"; 
      when 6456 => DO <= x"00000000"; 
      when 6457 => DO <= x"00000000"; 
      when 6458 => DO <= x"00000000"; 
      when 6459 => DO <= x"00000000"; 
      when 6460 => DO <= x"00000000"; 
      when 6461 => DO <= x"00000000"; 
      when 6462 => DO <= x"00000000"; 
      when 6463 => DO <= x"00000000"; 
      when 6464 => DO <= x"00000000"; 
      when 6465 => DO <= x"00000000"; 
      when 6466 => DO <= x"00000000"; 
      when 6467 => DO <= x"00000000"; 
      when 6468 => DO <= x"00000000"; 
      when 6469 => DO <= x"00000000"; 
      when 6470 => DO <= x"00000000"; 
      when 6471 => DO <= x"00000000"; 
      when 6472 => DO <= x"00000000"; 
      when 6473 => DO <= x"00000000"; 
      when 6474 => DO <= x"00000000"; 
      when 6475 => DO <= x"00000000"; 
      when 6476 => DO <= x"00000000"; 
      when 6477 => DO <= x"00000000"; 
      when 6478 => DO <= x"00000000"; 
      when 6479 => DO <= x"00000000"; 
      when 6480 => DO <= x"00000000"; 
      when 6481 => DO <= x"00000000"; 
      when 6482 => DO <= x"00000000"; 
      when 6483 => DO <= x"00000000"; 
      when 6484 => DO <= x"00000000"; 
      when 6485 => DO <= x"00000000"; 
      when 6486 => DO <= x"00000000"; 
      when 6487 => DO <= x"00000000"; 
      when 6488 => DO <= x"00000000"; 
      when 6489 => DO <= x"00000000"; 
      when 6490 => DO <= x"00000000"; 
      when 6491 => DO <= x"00000000"; 
      when 6492 => DO <= x"00000000"; 
      when 6493 => DO <= x"00000000"; 
      when 6494 => DO <= x"00000000"; 
      when 6495 => DO <= x"00000000"; 
      when 6496 => DO <= x"00000000"; 
      when 6497 => DO <= x"00000000"; 
      when 6498 => DO <= x"00000000"; 
      when 6499 => DO <= x"00000000"; 
      when 6500 => DO <= x"00000000"; 
      when 6501 => DO <= x"00000000"; 
      when 6502 => DO <= x"00000000"; 
      when 6503 => DO <= x"00000000"; 
      when 6504 => DO <= x"00000000"; 
      when 6505 => DO <= x"00000000"; 
      when 6506 => DO <= x"00000000"; 
      when 6507 => DO <= x"00000000"; 
      when 6508 => DO <= x"00000000"; 
      when 6509 => DO <= x"00000000"; 
      when 6510 => DO <= x"00000000"; 
      when 6511 => DO <= x"00000000"; 
      when 6512 => DO <= x"00000000"; 
      when 6513 => DO <= x"00000000"; 
      when 6514 => DO <= x"00000000"; 
      when 6515 => DO <= x"00000000"; 
      when 6516 => DO <= x"00000000"; 
      when 6517 => DO <= x"00000000"; 
      when 6518 => DO <= x"00000000"; 
      when 6519 => DO <= x"00000000"; 
      when 6520 => DO <= x"00000000"; 
      when 6521 => DO <= x"00000000"; 
      when 6522 => DO <= x"00000000"; 
      when 6523 => DO <= x"00000000"; 
      when 6524 => DO <= x"00000000"; 
      when 6525 => DO <= x"00000000"; 
      when 6526 => DO <= x"00000000"; 
      when 6527 => DO <= x"00000000"; 
      when 6528 => DO <= x"00000000"; 
      when 6529 => DO <= x"00000000"; 
      when 6530 => DO <= x"00000000"; 
      when 6531 => DO <= x"00000000"; 
      when 6532 => DO <= x"00000000"; 
      when 6533 => DO <= x"00000000"; 
      when 6534 => DO <= x"00000000"; 
      when 6535 => DO <= x"00000000"; 
      when 6536 => DO <= x"00000000"; 
      when 6537 => DO <= x"00000000"; 
      when 6538 => DO <= x"00000000"; 
      when 6539 => DO <= x"00000000"; 
      when 6540 => DO <= x"00000000"; 
      when 6541 => DO <= x"00000000"; 
      when 6542 => DO <= x"00000000"; 
      when 6543 => DO <= x"00000000"; 
      when 6544 => DO <= x"00000000"; 
      when 6545 => DO <= x"00000000"; 
      when 6546 => DO <= x"00000000"; 
      when 6547 => DO <= x"00000000"; 
      when 6548 => DO <= x"00000000"; 
      when 6549 => DO <= x"00000000"; 
      when 6550 => DO <= x"00000000"; 
      when 6551 => DO <= x"00000000"; 
      when 6552 => DO <= x"00000000"; 
      when 6553 => DO <= x"00000000"; 
      when 6554 => DO <= x"00000000"; 
      when 6555 => DO <= x"00000000"; 
      when 6556 => DO <= x"00000000"; 
      when 6557 => DO <= x"00000000"; 
      when 6558 => DO <= x"00000000"; 
      when 6559 => DO <= x"00000000"; 
      when 6560 => DO <= x"00000000"; 
      when 6561 => DO <= x"00000000"; 
      when 6562 => DO <= x"00000000"; 
      when 6563 => DO <= x"00000000"; 
      when 6564 => DO <= x"00000000"; 
      when 6565 => DO <= x"00000000"; 
      when 6566 => DO <= x"00000000"; 
      when 6567 => DO <= x"00000000"; 
      when 6568 => DO <= x"00000000"; 
      when 6569 => DO <= x"00000000"; 
      when 6570 => DO <= x"00000000"; 
      when 6571 => DO <= x"00000000"; 
      when 6572 => DO <= x"00000000"; 
      when 6573 => DO <= x"00000000"; 
      when 6574 => DO <= x"00000000"; 
      when 6575 => DO <= x"00000000"; 
      when 6576 => DO <= x"00000000"; 
      when 6577 => DO <= x"00000000"; 
      when 6578 => DO <= x"00000000"; 
      when 6579 => DO <= x"00000000"; 
      when 6580 => DO <= x"00000000"; 
      when 6581 => DO <= x"00000000"; 
      when 6582 => DO <= x"00000000"; 
      when 6583 => DO <= x"00000000"; 
      when 6584 => DO <= x"00000000"; 
      when 6585 => DO <= x"00000000"; 
      when 6586 => DO <= x"00000000"; 
      when 6587 => DO <= x"00000000"; 
      when 6588 => DO <= x"00000000"; 
      when 6589 => DO <= x"00000000"; 
      when 6590 => DO <= x"00000000"; 
      when 6591 => DO <= x"00000000"; 
      when 6592 => DO <= x"00000000"; 
      when 6593 => DO <= x"00000000"; 
      when 6594 => DO <= x"00000000"; 
      when 6595 => DO <= x"00000000"; 
      when 6596 => DO <= x"00000000"; 
      when 6597 => DO <= x"00000000"; 
      when 6598 => DO <= x"00000000"; 
      when 6599 => DO <= x"00000000"; 
      when 6600 => DO <= x"00000000"; 
      when 6601 => DO <= x"00000000"; 
      when 6602 => DO <= x"00000000"; 
      when 6603 => DO <= x"00000000"; 
      when 6604 => DO <= x"00000000"; 
      when 6605 => DO <= x"00000000"; 
      when 6606 => DO <= x"00000000"; 
      when 6607 => DO <= x"00000000"; 
      when 6608 => DO <= x"00000000"; 
      when 6609 => DO <= x"00000000"; 
      when 6610 => DO <= x"00000000"; 
      when 6611 => DO <= x"00000000"; 
      when 6612 => DO <= x"00000000"; 
      when 6613 => DO <= x"00000000"; 
      when 6614 => DO <= x"00000000"; 
      when 6615 => DO <= x"00000000"; 
      when 6616 => DO <= x"00000000"; 
      when 6617 => DO <= x"00000000"; 
      when 6618 => DO <= x"00000000"; 
      when 6619 => DO <= x"00000000"; 
      when 6620 => DO <= x"00000000"; 
      when 6621 => DO <= x"00000000"; 
      when 6622 => DO <= x"00000000"; 
      when 6623 => DO <= x"00000000"; 
      when 6624 => DO <= x"00000000"; 
      when 6625 => DO <= x"00000000"; 
      when 6626 => DO <= x"00000000"; 
      when 6627 => DO <= x"00000000"; 
      when 6628 => DO <= x"00000000"; 
      when 6629 => DO <= x"00000000"; 
      when 6630 => DO <= x"00000000"; 
      when 6631 => DO <= x"00000000"; 
      when 6632 => DO <= x"00000000"; 
      when 6633 => DO <= x"00000000"; 
      when 6634 => DO <= x"00000000"; 
      when 6635 => DO <= x"00000000"; 
      when 6636 => DO <= x"00000000"; 
      when 6637 => DO <= x"00000000"; 
      when 6638 => DO <= x"00000000"; 
      when 6639 => DO <= x"00000000"; 
      when 6640 => DO <= x"00000000"; 
      when 6641 => DO <= x"00000000"; 
      when 6642 => DO <= x"00000000"; 
      when 6643 => DO <= x"00000000"; 
      when 6644 => DO <= x"00000000"; 
      when 6645 => DO <= x"00000000"; 
      when 6646 => DO <= x"00000000"; 
      when 6647 => DO <= x"00000000"; 
      when 6648 => DO <= x"00000000"; 
      when 6649 => DO <= x"00000000"; 
      when 6650 => DO <= x"00000000"; 
      when 6651 => DO <= x"00000000"; 
      when 6652 => DO <= x"00000000"; 
      when 6653 => DO <= x"00000000"; 
      when 6654 => DO <= x"00000000"; 
      when 6655 => DO <= x"00000000"; 
      when 6656 => DO <= x"00000000"; 
      when 6657 => DO <= x"00000000"; 
      when 6658 => DO <= x"00000000"; 
      when 6659 => DO <= x"00000000"; 
      when 6660 => DO <= x"00000000"; 
      when 6661 => DO <= x"00000000"; 
      when 6662 => DO <= x"00000000"; 
      when 6663 => DO <= x"00000000"; 
      when 6664 => DO <= x"00000000"; 
      when 6665 => DO <= x"00000000"; 
      when 6666 => DO <= x"00000000"; 
      when 6667 => DO <= x"00000000"; 
      when 6668 => DO <= x"00000000"; 
      when 6669 => DO <= x"00000000"; 
      when 6670 => DO <= x"00000000"; 
      when 6671 => DO <= x"00000000"; 
      when 6672 => DO <= x"00000000"; 
      when 6673 => DO <= x"00000000"; 
      when 6674 => DO <= x"00000000"; 
      when 6675 => DO <= x"00000000"; 
      when 6676 => DO <= x"00000000"; 
      when 6677 => DO <= x"00000000"; 
      when 6678 => DO <= x"00000000"; 
      when 6679 => DO <= x"00000000"; 
      when 6680 => DO <= x"00000000"; 
      when 6681 => DO <= x"00000000"; 
      when 6682 => DO <= x"00000000"; 
      when 6683 => DO <= x"00000000"; 
      when 6684 => DO <= x"00000000"; 
      when 6685 => DO <= x"00000000"; 
      when 6686 => DO <= x"00000000"; 
      when 6687 => DO <= x"00000000"; 
      when 6688 => DO <= x"00000000"; 
      when 6689 => DO <= x"00000000"; 
      when 6690 => DO <= x"00000000"; 
      when 6691 => DO <= x"00000000"; 
      when 6692 => DO <= x"00000000"; 
      when 6693 => DO <= x"00000000"; 
      when 6694 => DO <= x"00000000"; 
      when 6695 => DO <= x"00000000"; 
      when 6696 => DO <= x"00000000"; 
      when 6697 => DO <= x"00000000"; 
      when 6698 => DO <= x"00000000"; 
      when 6699 => DO <= x"00000000"; 
      when 6700 => DO <= x"00000000"; 
      when 6701 => DO <= x"00000000"; 
      when 6702 => DO <= x"00000000"; 
      when 6703 => DO <= x"00000000"; 
      when 6704 => DO <= x"00000000"; 
      when 6705 => DO <= x"00000000"; 
      when 6706 => DO <= x"00000000"; 
      when 6707 => DO <= x"00000000"; 
      when 6708 => DO <= x"00000000"; 
      when 6709 => DO <= x"00000000"; 
      when 6710 => DO <= x"00000000"; 
      when 6711 => DO <= x"00000000"; 
      when 6712 => DO <= x"00000000"; 
      when 6713 => DO <= x"00000000"; 
      when 6714 => DO <= x"00000000"; 
      when 6715 => DO <= x"00000000"; 
      when 6716 => DO <= x"00000000"; 
      when 6717 => DO <= x"00000000"; 
      when 6718 => DO <= x"00000000"; 
      when 6719 => DO <= x"00000000"; 
      when 6720 => DO <= x"00000000"; 
      when 6721 => DO <= x"00000000"; 
      when 6722 => DO <= x"00000000"; 
      when 6723 => DO <= x"00000000"; 
      when 6724 => DO <= x"00000000"; 
      when 6725 => DO <= x"00000000"; 
      when 6726 => DO <= x"00000000"; 
      when 6727 => DO <= x"00000000"; 
      when 6728 => DO <= x"00000000"; 
      when 6729 => DO <= x"00000000"; 
      when 6730 => DO <= x"00000000"; 
      when 6731 => DO <= x"00000000"; 
      when 6732 => DO <= x"00000000"; 
      when 6733 => DO <= x"00000000"; 
      when 6734 => DO <= x"00000000"; 
      when 6735 => DO <= x"00000000"; 
      when 6736 => DO <= x"00000000"; 
      when 6737 => DO <= x"00000000"; 
      when 6738 => DO <= x"00000000"; 
      when 6739 => DO <= x"00000000"; 
      when 6740 => DO <= x"00000000"; 
      when 6741 => DO <= x"00000000"; 
      when 6742 => DO <= x"00000000"; 
      when 6743 => DO <= x"00000000"; 
      when 6744 => DO <= x"00000000"; 
      when 6745 => DO <= x"00000000"; 
      when 6746 => DO <= x"00000000"; 
      when 6747 => DO <= x"00000000"; 
      when 6748 => DO <= x"00000000"; 
      when 6749 => DO <= x"00000000"; 
      when 6750 => DO <= x"00000000"; 
      when 6751 => DO <= x"00000000"; 
      when 6752 => DO <= x"00000000"; 
      when 6753 => DO <= x"00000000"; 
      when 6754 => DO <= x"00000000"; 
      when 6755 => DO <= x"00000000"; 
      when 6756 => DO <= x"00000000"; 
      when 6757 => DO <= x"00000000"; 
      when 6758 => DO <= x"00000000"; 
      when 6759 => DO <= x"00000000"; 
      when 6760 => DO <= x"00000000"; 
      when 6761 => DO <= x"00000000"; 
      when 6762 => DO <= x"00000000"; 
      when 6763 => DO <= x"00000000"; 
      when 6764 => DO <= x"00000000"; 
      when 6765 => DO <= x"00000000"; 
      when 6766 => DO <= x"00000000"; 
      when 6767 => DO <= x"00000000"; 
      when 6768 => DO <= x"00000000"; 
      when 6769 => DO <= x"00000000"; 
      when 6770 => DO <= x"00000000"; 
      when 6771 => DO <= x"00000000"; 
      when 6772 => DO <= x"00000000"; 
      when 6773 => DO <= x"00000000"; 
      when 6774 => DO <= x"00000000"; 
      when 6775 => DO <= x"00000000"; 
      when 6776 => DO <= x"00000000"; 
      when 6777 => DO <= x"00000000"; 
      when 6778 => DO <= x"00000000"; 
      when 6779 => DO <= x"00000000"; 
      when 6780 => DO <= x"00000000"; 
      when 6781 => DO <= x"00000000"; 
      when 6782 => DO <= x"00000000"; 
      when 6783 => DO <= x"00000000"; 
      when 6784 => DO <= x"00000000"; 
      when 6785 => DO <= x"00000000"; 
      when 6786 => DO <= x"00000000"; 
      when 6787 => DO <= x"00000000"; 
      when 6788 => DO <= x"00000000"; 
      when 6789 => DO <= x"00000000"; 
      when 6790 => DO <= x"00000000"; 
      when 6791 => DO <= x"00000000"; 
      when 6792 => DO <= x"00000000"; 
      when 6793 => DO <= x"00000000"; 
      when 6794 => DO <= x"00000000"; 
      when 6795 => DO <= x"00000000"; 
      when 6796 => DO <= x"00000000"; 
      when 6797 => DO <= x"00000000"; 
      when 6798 => DO <= x"00000000"; 
      when 6799 => DO <= x"00000000"; 
      when 6800 => DO <= x"00000000"; 
      when 6801 => DO <= x"00000000"; 
      when 6802 => DO <= x"00000000"; 
      when 6803 => DO <= x"00000000"; 
      when 6804 => DO <= x"00000000"; 
      when 6805 => DO <= x"00000000"; 
      when 6806 => DO <= x"00000000"; 
      when 6807 => DO <= x"00000000"; 
      when 6808 => DO <= x"00000000"; 
      when 6809 => DO <= x"00000000"; 
      when 6810 => DO <= x"00000000"; 
      when 6811 => DO <= x"00000000"; 
      when 6812 => DO <= x"00000000"; 
      when 6813 => DO <= x"00000000"; 
      when 6814 => DO <= x"00000000"; 
      when 6815 => DO <= x"00000000"; 
      when 6816 => DO <= x"00000000"; 
      when 6817 => DO <= x"00000000"; 
      when 6818 => DO <= x"00000000"; 
      when 6819 => DO <= x"00000000"; 
      when 6820 => DO <= x"00000000"; 
      when 6821 => DO <= x"00000000"; 
      when 6822 => DO <= x"00000000"; 
      when 6823 => DO <= x"00000000"; 
      when 6824 => DO <= x"00000000"; 
      when 6825 => DO <= x"00000000"; 
      when 6826 => DO <= x"00000000"; 
      when 6827 => DO <= x"00000000"; 
      when 6828 => DO <= x"00000000"; 
      when 6829 => DO <= x"00000000"; 
      when 6830 => DO <= x"00000000"; 
      when 6831 => DO <= x"00000000"; 
      when 6832 => DO <= x"00000000"; 
      when 6833 => DO <= x"00000000"; 
      when 6834 => DO <= x"00000000"; 
      when 6835 => DO <= x"00000000"; 
      when 6836 => DO <= x"00000000"; 
      when 6837 => DO <= x"00000000"; 
      when 6838 => DO <= x"00000000"; 
      when 6839 => DO <= x"00000000"; 
      when 6840 => DO <= x"00000000"; 
      when 6841 => DO <= x"00000000"; 
      when 6842 => DO <= x"00000000"; 
      when 6843 => DO <= x"00000000"; 
      when 6844 => DO <= x"00000000"; 
      when 6845 => DO <= x"00000000"; 
      when 6846 => DO <= x"00000000"; 
      when 6847 => DO <= x"00000000"; 
      when 6848 => DO <= x"00000000"; 
      when 6849 => DO <= x"00000000"; 
      when 6850 => DO <= x"00000000"; 
      when 6851 => DO <= x"00000000"; 
      when 6852 => DO <= x"00000000"; 
      when 6853 => DO <= x"00000000"; 
      when 6854 => DO <= x"00000000"; 
      when 6855 => DO <= x"00000000"; 
      when 6856 => DO <= x"00000000"; 
      when 6857 => DO <= x"00000000"; 
      when 6858 => DO <= x"00000000"; 
      when 6859 => DO <= x"00000000"; 
      when 6860 => DO <= x"00000000"; 
      when 6861 => DO <= x"00000000"; 
      when 6862 => DO <= x"00000000"; 
      when 6863 => DO <= x"00000000"; 
      when 6864 => DO <= x"00000000"; 
      when 6865 => DO <= x"00000000"; 
      when 6866 => DO <= x"00000000"; 
      when 6867 => DO <= x"00000000"; 
      when 6868 => DO <= x"00000000"; 
      when 6869 => DO <= x"00000000"; 
      when 6870 => DO <= x"00000000"; 
      when 6871 => DO <= x"00000000"; 
      when 6872 => DO <= x"00000000"; 
      when 6873 => DO <= x"00000000"; 
      when 6874 => DO <= x"00000000"; 
      when 6875 => DO <= x"00000000"; 
      when 6876 => DO <= x"00000000"; 
      when 6877 => DO <= x"00000000"; 
      when 6878 => DO <= x"00000000"; 
      when 6879 => DO <= x"00000000"; 
      when 6880 => DO <= x"00000000"; 
      when 6881 => DO <= x"00000000"; 
      when 6882 => DO <= x"00000000"; 
      when 6883 => DO <= x"00000000"; 
      when 6884 => DO <= x"00000000"; 
      when 6885 => DO <= x"00000000"; 
      when 6886 => DO <= x"00000000"; 
      when 6887 => DO <= x"00000000"; 
      when 6888 => DO <= x"00000000"; 
      when 6889 => DO <= x"00000000"; 
      when 6890 => DO <= x"00000000"; 
      when 6891 => DO <= x"00000000"; 
      when 6892 => DO <= x"00000000"; 
      when 6893 => DO <= x"00000000"; 
      when 6894 => DO <= x"00000000"; 
      when 6895 => DO <= x"00000000"; 
      when 6896 => DO <= x"00000000"; 
      when 6897 => DO <= x"00000000"; 
      when 6898 => DO <= x"00000000"; 
      when 6899 => DO <= x"00000000"; 
      when 6900 => DO <= x"00000000"; 
      when 6901 => DO <= x"00000000"; 
      when 6902 => DO <= x"00000000"; 
      when 6903 => DO <= x"00000000"; 
      when 6904 => DO <= x"00000000"; 
      when 6905 => DO <= x"00000000"; 
      when 6906 => DO <= x"00000000"; 
      when 6907 => DO <= x"00000000"; 
      when 6908 => DO <= x"00000000"; 
      when 6909 => DO <= x"00000000"; 
      when 6910 => DO <= x"00000000"; 
      when 6911 => DO <= x"00000000"; 
      when 6912 => DO <= x"00000000"; 
      when 6913 => DO <= x"00000000"; 
      when 6914 => DO <= x"00000000"; 
      when 6915 => DO <= x"00000000"; 
      when 6916 => DO <= x"00000000"; 
      when 6917 => DO <= x"00000000"; 
      when 6918 => DO <= x"00000000"; 
      when 6919 => DO <= x"00000000"; 
      when 6920 => DO <= x"00000000"; 
      when 6921 => DO <= x"00000000"; 
      when 6922 => DO <= x"00000000"; 
      when 6923 => DO <= x"00000000"; 
      when 6924 => DO <= x"00000000"; 
      when 6925 => DO <= x"00000000"; 
      when 6926 => DO <= x"00000000"; 
      when 6927 => DO <= x"00000000"; 
      when 6928 => DO <= x"00000000"; 
      when 6929 => DO <= x"00000000"; 
      when 6930 => DO <= x"00000000"; 
      when 6931 => DO <= x"00000000"; 
      when 6932 => DO <= x"00000000"; 
      when 6933 => DO <= x"00000000"; 
      when 6934 => DO <= x"00000000"; 
      when 6935 => DO <= x"00000000"; 
      when 6936 => DO <= x"00000000"; 
      when 6937 => DO <= x"00000000"; 
      when 6938 => DO <= x"00000000"; 
      when 6939 => DO <= x"00000000"; 
      when 6940 => DO <= x"00000000"; 
      when 6941 => DO <= x"00000000"; 
      when 6942 => DO <= x"00000000"; 
      when 6943 => DO <= x"00000000"; 
      when 6944 => DO <= x"00000000"; 
      when 6945 => DO <= x"00000000"; 
      when 6946 => DO <= x"00000000"; 
      when 6947 => DO <= x"00000000"; 
      when 6948 => DO <= x"00000000"; 
      when 6949 => DO <= x"00000000"; 
      when 6950 => DO <= x"00000000"; 
      when 6951 => DO <= x"00000000"; 
      when 6952 => DO <= x"00000000"; 
      when 6953 => DO <= x"00000000"; 
      when 6954 => DO <= x"00000000"; 
      when 6955 => DO <= x"00000000"; 
      when 6956 => DO <= x"00000000"; 
      when 6957 => DO <= x"00000000"; 
      when 6958 => DO <= x"00000000"; 
      when 6959 => DO <= x"00000000"; 
      when 6960 => DO <= x"00000000"; 
      when 6961 => DO <= x"00000000"; 
      when 6962 => DO <= x"00000000"; 
      when 6963 => DO <= x"00000000"; 
      when 6964 => DO <= x"00000000"; 
      when 6965 => DO <= x"00000000"; 
      when 6966 => DO <= x"00000000"; 
      when 6967 => DO <= x"00000000"; 
      when 6968 => DO <= x"00000000"; 
      when 6969 => DO <= x"00000000"; 
      when 6970 => DO <= x"00000000"; 
      when 6971 => DO <= x"00000000"; 
      when 6972 => DO <= x"00000000"; 
      when 6973 => DO <= x"00000000"; 
      when 6974 => DO <= x"00000000"; 
      when 6975 => DO <= x"00000000"; 
      when 6976 => DO <= x"00000000"; 
      when 6977 => DO <= x"00000000"; 
      when 6978 => DO <= x"00000000"; 
      when 6979 => DO <= x"00000000"; 
      when 6980 => DO <= x"00000000"; 
      when 6981 => DO <= x"00000000"; 
      when 6982 => DO <= x"00000000"; 
      when 6983 => DO <= x"00000000"; 
      when 6984 => DO <= x"00000000"; 
      when 6985 => DO <= x"00000000"; 
      when 6986 => DO <= x"00000000"; 
      when 6987 => DO <= x"00000000"; 
      when 6988 => DO <= x"00000000"; 
      when 6989 => DO <= x"00000000"; 
      when 6990 => DO <= x"00000000"; 
      when 6991 => DO <= x"00000000"; 
      when 6992 => DO <= x"00000000"; 
      when 6993 => DO <= x"00000000"; 
      when 6994 => DO <= x"00000000"; 
      when 6995 => DO <= x"00000000"; 
      when 6996 => DO <= x"00000000"; 
      when 6997 => DO <= x"00000000"; 
      when 6998 => DO <= x"00000000"; 
      when 6999 => DO <= x"00000000"; 
      when 7000 => DO <= x"00000000"; 
      when 7001 => DO <= x"00000000"; 
      when 7002 => DO <= x"00000000"; 
      when 7003 => DO <= x"00000000"; 
      when 7004 => DO <= x"00000000"; 
      when 7005 => DO <= x"00000000"; 
      when 7006 => DO <= x"00000000"; 
      when 7007 => DO <= x"00000000"; 
      when 7008 => DO <= x"00000000"; 
      when 7009 => DO <= x"00000000"; 
      when 7010 => DO <= x"00000000"; 
      when 7011 => DO <= x"00000000"; 
      when 7012 => DO <= x"00000000"; 
      when 7013 => DO <= x"00000000"; 
      when 7014 => DO <= x"00000000"; 
      when 7015 => DO <= x"00000000"; 
      when 7016 => DO <= x"00000000"; 
      when 7017 => DO <= x"00000000"; 
      when 7018 => DO <= x"00000000"; 
      when 7019 => DO <= x"00000000"; 
      when 7020 => DO <= x"00000000"; 
      when 7021 => DO <= x"00000000"; 
      when 7022 => DO <= x"00000000"; 
      when 7023 => DO <= x"00000000"; 
      when 7024 => DO <= x"00000000"; 
      when 7025 => DO <= x"00000000"; 
      when 7026 => DO <= x"00000000"; 
      when 7027 => DO <= x"00000000"; 
      when 7028 => DO <= x"00000000"; 
      when 7029 => DO <= x"00000000"; 
      when 7030 => DO <= x"00000000"; 
      when 7031 => DO <= x"00000000"; 
      when 7032 => DO <= x"00000000"; 
      when 7033 => DO <= x"00000000"; 
      when 7034 => DO <= x"00000000"; 
      when 7035 => DO <= x"00000000"; 
      when 7036 => DO <= x"00000000"; 
      when 7037 => DO <= x"00000000"; 
      when 7038 => DO <= x"00000000"; 
      when 7039 => DO <= x"00000000"; 
      when 7040 => DO <= x"00000000"; 
      when 7041 => DO <= x"00000000"; 
      when 7042 => DO <= x"00000000"; 
      when 7043 => DO <= x"00000000"; 
      when 7044 => DO <= x"00000000"; 
      when 7045 => DO <= x"00000000"; 
      when 7046 => DO <= x"00000000"; 
      when 7047 => DO <= x"00000000"; 
      when 7048 => DO <= x"00000000"; 
      when 7049 => DO <= x"00000000"; 
      when 7050 => DO <= x"00000000"; 
      when 7051 => DO <= x"00000000"; 
      when 7052 => DO <= x"00000000"; 
      when 7053 => DO <= x"00000000"; 
      when 7054 => DO <= x"00000000"; 
      when 7055 => DO <= x"00000000"; 
      when 7056 => DO <= x"00000000"; 
      when 7057 => DO <= x"00000000"; 
      when 7058 => DO <= x"00000000"; 
      when 7059 => DO <= x"00000000"; 
      when 7060 => DO <= x"00000000"; 
      when 7061 => DO <= x"00000000"; 
      when 7062 => DO <= x"00000000"; 
      when 7063 => DO <= x"00000000"; 
      when 7064 => DO <= x"00000000"; 
      when 7065 => DO <= x"00000000"; 
      when 7066 => DO <= x"00000000"; 
      when 7067 => DO <= x"00000000"; 
      when 7068 => DO <= x"00000000"; 
      when 7069 => DO <= x"00000000"; 
      when 7070 => DO <= x"00000000"; 
      when 7071 => DO <= x"00000000"; 
      when 7072 => DO <= x"00000000"; 
      when 7073 => DO <= x"00000000"; 
      when 7074 => DO <= x"00000000"; 
      when 7075 => DO <= x"00000000"; 
      when 7076 => DO <= x"00000000"; 
      when 7077 => DO <= x"00000000"; 
      when 7078 => DO <= x"00000000"; 
      when 7079 => DO <= x"00000000"; 
      when 7080 => DO <= x"00000000"; 
      when 7081 => DO <= x"00000000"; 
      when 7082 => DO <= x"00000000"; 
      when 7083 => DO <= x"00000000"; 
      when 7084 => DO <= x"00000000"; 
      when 7085 => DO <= x"00000000"; 
      when 7086 => DO <= x"00000000"; 
      when 7087 => DO <= x"00000000"; 
      when 7088 => DO <= x"00000000"; 
      when 7089 => DO <= x"00000000"; 
      when 7090 => DO <= x"00000000"; 
      when 7091 => DO <= x"00000000"; 
      when 7092 => DO <= x"00000000"; 
      when 7093 => DO <= x"00000000"; 
      when 7094 => DO <= x"00000000"; 
      when 7095 => DO <= x"00000000"; 
      when 7096 => DO <= x"00000000"; 
      when 7097 => DO <= x"00000000"; 
      when 7098 => DO <= x"00000000"; 
      when 7099 => DO <= x"00000000"; 
      when 7100 => DO <= x"00000000"; 
      when 7101 => DO <= x"00000000"; 
      when 7102 => DO <= x"00000000"; 
      when 7103 => DO <= x"00000000"; 
      when 7104 => DO <= x"00000000"; 
      when 7105 => DO <= x"00000000"; 
      when 7106 => DO <= x"00000000"; 
      when 7107 => DO <= x"00000000"; 
      when 7108 => DO <= x"00000000"; 
      when 7109 => DO <= x"00000000"; 
      when 7110 => DO <= x"00000000"; 
      when 7111 => DO <= x"00000000"; 
      when 7112 => DO <= x"00000000"; 
      when 7113 => DO <= x"00000000"; 
      when 7114 => DO <= x"00000000"; 
      when 7115 => DO <= x"00000000"; 
      when 7116 => DO <= x"00000000"; 
      when 7117 => DO <= x"00000000"; 
      when 7118 => DO <= x"00000000"; 
      when 7119 => DO <= x"00000000"; 
      when 7120 => DO <= x"00000000"; 
      when 7121 => DO <= x"00000000"; 
      when 7122 => DO <= x"00000000"; 
      when 7123 => DO <= x"00000000"; 
      when 7124 => DO <= x"00000000"; 
      when 7125 => DO <= x"00000000"; 
      when 7126 => DO <= x"00000000"; 
      when 7127 => DO <= x"00000000"; 
      when 7128 => DO <= x"00000000"; 
      when 7129 => DO <= x"00000000"; 
      when 7130 => DO <= x"00000000"; 
      when 7131 => DO <= x"00000000"; 
      when 7132 => DO <= x"00000000"; 
      when 7133 => DO <= x"00000000"; 
      when 7134 => DO <= x"00000000"; 
      when 7135 => DO <= x"00000000"; 
      when 7136 => DO <= x"00000000"; 
      when 7137 => DO <= x"00000000"; 
      when 7138 => DO <= x"00000000"; 
      when 7139 => DO <= x"00000000"; 
      when 7140 => DO <= x"00000000"; 
      when 7141 => DO <= x"00000000"; 
      when 7142 => DO <= x"00000000"; 
      when 7143 => DO <= x"00000000"; 
      when 7144 => DO <= x"00000000"; 
      when 7145 => DO <= x"00000000"; 
      when 7146 => DO <= x"00000000"; 
      when 7147 => DO <= x"00000000"; 
      when 7148 => DO <= x"00000000"; 
      when 7149 => DO <= x"00000000"; 
      when 7150 => DO <= x"00000000"; 
      when 7151 => DO <= x"00000000"; 
      when 7152 => DO <= x"00000000"; 
      when 7153 => DO <= x"00000000"; 
      when 7154 => DO <= x"00000000"; 
      when 7155 => DO <= x"00000000"; 
      when 7156 => DO <= x"00000000"; 
      when 7157 => DO <= x"00000000"; 
      when 7158 => DO <= x"00000000"; 
      when 7159 => DO <= x"00000000"; 
      when 7160 => DO <= x"00000000"; 
      when 7161 => DO <= x"00000000"; 
      when 7162 => DO <= x"00000000"; 
      when 7163 => DO <= x"00000000"; 
      when 7164 => DO <= x"00000000"; 
      when 7165 => DO <= x"00000000"; 
      when 7166 => DO <= x"00000000"; 
      when 7167 => DO <= x"00000000"; 
      when 7168 => DO <= x"00000000"; 
      when 7169 => DO <= x"00000000"; 
      when 7170 => DO <= x"00000000"; 
      when 7171 => DO <= x"00000000"; 
      when 7172 => DO <= x"00000000"; 
      when 7173 => DO <= x"00000000"; 
      when 7174 => DO <= x"00000000"; 
      when 7175 => DO <= x"00000000"; 
      when 7176 => DO <= x"00000000"; 
      when 7177 => DO <= x"00000000"; 
      when 7178 => DO <= x"00000000"; 
      when 7179 => DO <= x"00000000"; 
      when 7180 => DO <= x"00000000"; 
      when 7181 => DO <= x"00000000"; 
      when 7182 => DO <= x"00000000"; 
      when 7183 => DO <= x"00000000"; 
      when 7184 => DO <= x"00000000"; 
      when 7185 => DO <= x"00000000"; 
      when 7186 => DO <= x"00000000"; 
      when 7187 => DO <= x"00000000"; 
      when 7188 => DO <= x"00000000"; 
      when 7189 => DO <= x"00000000"; 
      when 7190 => DO <= x"00000000"; 
      when 7191 => DO <= x"00000000"; 
      when 7192 => DO <= x"00000000"; 
      when 7193 => DO <= x"00000000"; 
      when 7194 => DO <= x"00000000"; 
      when 7195 => DO <= x"00000000"; 
      when 7196 => DO <= x"00000000"; 
      when 7197 => DO <= x"00000000"; 
      when 7198 => DO <= x"00000000"; 
      when 7199 => DO <= x"00000000"; 
      when 7200 => DO <= x"00000000"; 
      when 7201 => DO <= x"00000000"; 
      when 7202 => DO <= x"00000000"; 
      when 7203 => DO <= x"00000000"; 
      when 7204 => DO <= x"00000000"; 
      when 7205 => DO <= x"00000000"; 
      when 7206 => DO <= x"00000000"; 
      when 7207 => DO <= x"00000000"; 
      when 7208 => DO <= x"00000000"; 
      when 7209 => DO <= x"00000000"; 
      when 7210 => DO <= x"00000000"; 
      when 7211 => DO <= x"00000000"; 
      when 7212 => DO <= x"00000000"; 
      when 7213 => DO <= x"00000000"; 
      when 7214 => DO <= x"00000000"; 
      when 7215 => DO <= x"00000000"; 
      when 7216 => DO <= x"00000000"; 
      when 7217 => DO <= x"00000000"; 
      when 7218 => DO <= x"00000000"; 
      when 7219 => DO <= x"00000000"; 
      when 7220 => DO <= x"00000000"; 
      when 7221 => DO <= x"00000000"; 
      when 7222 => DO <= x"00000000"; 
      when 7223 => DO <= x"00000000"; 
      when 7224 => DO <= x"00000000"; 
      when 7225 => DO <= x"00000000"; 
      when 7226 => DO <= x"00000000"; 
      when 7227 => DO <= x"00000000"; 
      when 7228 => DO <= x"00000000"; 
      when 7229 => DO <= x"00000000"; 
      when 7230 => DO <= x"00000000"; 
      when 7231 => DO <= x"00000000"; 
      when 7232 => DO <= x"00000000"; 
      when 7233 => DO <= x"00000000"; 
      when 7234 => DO <= x"00000000"; 
      when 7235 => DO <= x"00000000"; 
      when 7236 => DO <= x"00000000"; 
      when 7237 => DO <= x"00000000"; 
      when 7238 => DO <= x"00000000"; 
      when 7239 => DO <= x"00000000"; 
      when 7240 => DO <= x"00000000"; 
      when 7241 => DO <= x"00000000"; 
      when 7242 => DO <= x"00000000"; 
      when 7243 => DO <= x"00000000"; 
      when 7244 => DO <= x"00000000"; 
      when 7245 => DO <= x"00000000"; 
      when 7246 => DO <= x"00000000"; 
      when 7247 => DO <= x"00000000"; 
      when 7248 => DO <= x"00000000"; 
      when 7249 => DO <= x"00000000"; 
      when 7250 => DO <= x"00000000"; 
      when 7251 => DO <= x"00000000"; 
      when 7252 => DO <= x"00000000"; 
      when 7253 => DO <= x"00000000"; 
      when 7254 => DO <= x"00000000"; 
      when 7255 => DO <= x"00000000"; 
      when 7256 => DO <= x"00000000"; 
      when 7257 => DO <= x"00000000"; 
      when 7258 => DO <= x"00000000"; 
      when 7259 => DO <= x"00000000"; 
      when 7260 => DO <= x"00000000"; 
      when 7261 => DO <= x"00000000"; 
      when 7262 => DO <= x"00000000"; 
      when 7263 => DO <= x"00000000"; 
      when 7264 => DO <= x"00000000"; 
      when 7265 => DO <= x"00000000"; 
      when 7266 => DO <= x"00000000"; 
      when 7267 => DO <= x"00000000"; 
      when 7268 => DO <= x"00000000"; 
      when 7269 => DO <= x"00000000"; 
      when 7270 => DO <= x"00000000"; 
      when 7271 => DO <= x"00000000"; 
      when 7272 => DO <= x"00000000"; 
      when 7273 => DO <= x"00000000"; 
      when 7274 => DO <= x"00000000"; 
      when 7275 => DO <= x"00000000"; 
      when 7276 => DO <= x"00000000"; 
      when 7277 => DO <= x"00000000"; 
      when 7278 => DO <= x"00000000"; 
      when 7279 => DO <= x"00000000"; 
      when 7280 => DO <= x"00000000"; 
      when 7281 => DO <= x"00000000"; 
      when 7282 => DO <= x"00000000"; 
      when 7283 => DO <= x"00000000"; 
      when 7284 => DO <= x"00000000"; 
      when 7285 => DO <= x"00000000"; 
      when 7286 => DO <= x"00000000"; 
      when 7287 => DO <= x"00000000"; 
      when 7288 => DO <= x"00000000"; 
      when 7289 => DO <= x"00000000"; 
      when 7290 => DO <= x"00000000"; 
      when 7291 => DO <= x"00000000"; 
      when 7292 => DO <= x"00000000"; 
      when 7293 => DO <= x"00000000"; 
      when 7294 => DO <= x"00000000"; 
      when 7295 => DO <= x"00000000"; 
      when 7296 => DO <= x"00000000"; 
      when 7297 => DO <= x"00000000"; 
      when 7298 => DO <= x"00000000"; 
      when 7299 => DO <= x"00000000"; 
      when 7300 => DO <= x"00000000"; 
      when 7301 => DO <= x"00000000"; 
      when 7302 => DO <= x"00000000"; 
      when 7303 => DO <= x"00000000"; 
      when 7304 => DO <= x"00000000"; 
      when 7305 => DO <= x"00000000"; 
      when 7306 => DO <= x"00000000"; 
      when 7307 => DO <= x"00000000"; 
      when 7308 => DO <= x"00000000"; 
      when 7309 => DO <= x"00000000"; 
      when 7310 => DO <= x"00000000"; 
      when 7311 => DO <= x"00000000"; 
      when 7312 => DO <= x"00000000"; 
      when 7313 => DO <= x"00000000"; 
      when 7314 => DO <= x"00000000"; 
      when 7315 => DO <= x"00000000"; 
      when 7316 => DO <= x"00000000"; 
      when 7317 => DO <= x"00000000"; 
      when 7318 => DO <= x"00000000"; 
      when 7319 => DO <= x"00000000"; 
      when 7320 => DO <= x"00000000"; 
      when 7321 => DO <= x"00000000"; 
      when 7322 => DO <= x"00000000"; 
      when 7323 => DO <= x"00000000"; 
      when 7324 => DO <= x"00000000"; 
      when 7325 => DO <= x"00000000"; 
      when 7326 => DO <= x"00000000"; 
      when 7327 => DO <= x"00000000"; 
      when 7328 => DO <= x"00000000"; 
      when 7329 => DO <= x"00000000"; 
      when 7330 => DO <= x"00000000"; 
      when 7331 => DO <= x"00000000"; 
      when 7332 => DO <= x"00000000"; 
      when 7333 => DO <= x"00000000"; 
      when 7334 => DO <= x"00000000"; 
      when 7335 => DO <= x"00000000"; 
      when 7336 => DO <= x"00000000"; 
      when 7337 => DO <= x"00000000"; 
      when 7338 => DO <= x"00000000"; 
      when 7339 => DO <= x"00000000"; 
      when 7340 => DO <= x"00000000"; 
      when 7341 => DO <= x"00000000"; 
      when 7342 => DO <= x"00000000"; 
      when 7343 => DO <= x"00000000"; 
      when 7344 => DO <= x"00000000"; 
      when 7345 => DO <= x"00000000"; 
      when 7346 => DO <= x"00000000"; 
      when 7347 => DO <= x"00000000"; 
      when 7348 => DO <= x"00000000"; 
      when 7349 => DO <= x"00000000"; 
      when 7350 => DO <= x"00000000"; 
      when 7351 => DO <= x"00000000"; 
      when 7352 => DO <= x"00000000"; 
      when 7353 => DO <= x"00000000"; 
      when 7354 => DO <= x"00000000"; 
      when 7355 => DO <= x"00000000"; 
      when 7356 => DO <= x"00000000"; 
      when 7357 => DO <= x"00000000"; 
      when 7358 => DO <= x"00000000"; 
      when 7359 => DO <= x"00000000"; 
      when 7360 => DO <= x"00000000"; 
      when 7361 => DO <= x"00000000"; 
      when 7362 => DO <= x"00000000"; 
      when 7363 => DO <= x"00000000"; 
      when 7364 => DO <= x"00000000"; 
      when 7365 => DO <= x"00000000"; 
      when 7366 => DO <= x"00000000"; 
      when 7367 => DO <= x"00000000"; 
      when 7368 => DO <= x"00000000"; 
      when 7369 => DO <= x"00000000"; 
      when 7370 => DO <= x"00000000"; 
      when 7371 => DO <= x"00000000"; 
      when 7372 => DO <= x"00000000"; 
      when 7373 => DO <= x"00000000"; 
      when 7374 => DO <= x"00000000"; 
      when 7375 => DO <= x"00000000"; 
      when 7376 => DO <= x"00000000"; 
      when 7377 => DO <= x"00000000"; 
      when 7378 => DO <= x"00000000"; 
      when 7379 => DO <= x"00000000"; 
      when 7380 => DO <= x"00000000"; 
      when 7381 => DO <= x"00000000"; 
      when 7382 => DO <= x"00000000"; 
      when 7383 => DO <= x"00000000"; 
      when 7384 => DO <= x"00000000"; 
      when 7385 => DO <= x"00000000"; 
      when 7386 => DO <= x"00000000"; 
      when 7387 => DO <= x"00000000"; 
      when 7388 => DO <= x"00000000"; 
      when 7389 => DO <= x"00000000"; 
      when 7390 => DO <= x"00000000"; 
      when 7391 => DO <= x"00000000"; 
      when 7392 => DO <= x"00000000"; 
      when 7393 => DO <= x"00000000"; 
      when 7394 => DO <= x"00000000"; 
      when 7395 => DO <= x"00000000"; 
      when 7396 => DO <= x"00000000"; 
      when 7397 => DO <= x"00000000"; 
      when 7398 => DO <= x"00000000"; 
      when 7399 => DO <= x"00000000"; 
      when 7400 => DO <= x"00000000"; 
      when 7401 => DO <= x"00000000"; 
      when 7402 => DO <= x"00000000"; 
      when 7403 => DO <= x"00000000"; 
      when 7404 => DO <= x"00000000"; 
      when 7405 => DO <= x"00000000"; 
      when 7406 => DO <= x"00000000"; 
      when 7407 => DO <= x"00000000"; 
      when 7408 => DO <= x"00000000"; 
      when 7409 => DO <= x"00000000"; 
      when 7410 => DO <= x"00000000"; 
      when 7411 => DO <= x"00000000"; 
      when 7412 => DO <= x"00000000"; 
      when 7413 => DO <= x"00000000"; 
      when 7414 => DO <= x"00000000"; 
      when 7415 => DO <= x"00000000"; 
      when 7416 => DO <= x"00000000"; 
      when 7417 => DO <= x"00000000"; 
      when 7418 => DO <= x"00000000"; 
      when 7419 => DO <= x"00000000"; 
      when 7420 => DO <= x"00000000"; 
      when 7421 => DO <= x"00000000"; 
      when 7422 => DO <= x"00000000"; 
      when 7423 => DO <= x"00000000"; 
      when 7424 => DO <= x"00000000"; 
      when 7425 => DO <= x"00000000"; 
      when 7426 => DO <= x"00000000"; 
      when 7427 => DO <= x"00000000"; 
      when 7428 => DO <= x"00000000"; 
      when 7429 => DO <= x"00000000"; 
      when 7430 => DO <= x"00000000"; 
      when 7431 => DO <= x"00000000"; 
      when 7432 => DO <= x"00000000"; 
      when 7433 => DO <= x"00000000"; 
      when 7434 => DO <= x"00000000"; 
      when 7435 => DO <= x"00000000"; 
      when 7436 => DO <= x"00000000"; 
      when 7437 => DO <= x"00000000"; 
      when 7438 => DO <= x"00000000"; 
      when 7439 => DO <= x"00000000"; 
      when 7440 => DO <= x"00000000"; 
      when 7441 => DO <= x"00000000"; 
      when 7442 => DO <= x"00000000"; 
      when 7443 => DO <= x"00000000"; 
      when 7444 => DO <= x"00000000"; 
      when 7445 => DO <= x"00000000"; 
      when 7446 => DO <= x"00000000"; 
      when 7447 => DO <= x"00000000"; 
      when 7448 => DO <= x"00000000"; 
      when 7449 => DO <= x"00000000"; 
      when 7450 => DO <= x"00000000"; 
      when 7451 => DO <= x"00000000"; 
      when 7452 => DO <= x"00000000"; 
      when 7453 => DO <= x"00000000"; 
      when 7454 => DO <= x"00000000"; 
      when 7455 => DO <= x"00000000"; 
      when 7456 => DO <= x"00000000"; 
      when 7457 => DO <= x"00000000"; 
      when 7458 => DO <= x"00000000"; 
      when 7459 => DO <= x"00000000"; 
      when 7460 => DO <= x"00000000"; 
      when 7461 => DO <= x"00000000"; 
      when 7462 => DO <= x"00000000"; 
      when 7463 => DO <= x"00000000"; 
      when 7464 => DO <= x"00000000"; 
      when 7465 => DO <= x"00000000"; 
      when 7466 => DO <= x"00000000"; 
      when 7467 => DO <= x"00000000"; 
      when 7468 => DO <= x"00000000"; 
      when 7469 => DO <= x"00000000"; 
      when 7470 => DO <= x"00000000"; 
      when 7471 => DO <= x"00000000"; 
      when 7472 => DO <= x"00000000"; 
      when 7473 => DO <= x"00000000"; 
      when 7474 => DO <= x"00000000"; 
      when 7475 => DO <= x"00000000"; 
      when 7476 => DO <= x"00000000"; 
      when 7477 => DO <= x"00000000"; 
      when 7478 => DO <= x"00000000"; 
      when 7479 => DO <= x"00000000"; 
      when 7480 => DO <= x"00000000"; 
      when 7481 => DO <= x"00000000"; 
      when 7482 => DO <= x"00000000"; 
      when 7483 => DO <= x"00000000"; 
      when 7484 => DO <= x"00000000"; 
      when 7485 => DO <= x"00000000"; 
      when 7486 => DO <= x"00000000"; 
      when 7487 => DO <= x"00000000"; 
      when 7488 => DO <= x"00000000"; 
      when 7489 => DO <= x"00000000"; 
      when 7490 => DO <= x"00000000"; 
      when 7491 => DO <= x"00000000"; 
      when 7492 => DO <= x"00000000"; 
      when 7493 => DO <= x"00000000"; 
      when 7494 => DO <= x"00000000"; 
      when 7495 => DO <= x"00000000"; 
      when 7496 => DO <= x"00000000"; 
      when 7497 => DO <= x"00000000"; 
      when 7498 => DO <= x"00000000"; 
      when 7499 => DO <= x"00000000"; 
      when 7500 => DO <= x"00000000"; 
      when 7501 => DO <= x"00000000"; 
      when 7502 => DO <= x"00000000"; 
      when 7503 => DO <= x"00000000"; 
      when 7504 => DO <= x"00000000"; 
      when 7505 => DO <= x"00000000"; 
      when 7506 => DO <= x"00000000"; 
      when 7507 => DO <= x"00000000"; 
      when 7508 => DO <= x"00000000"; 
      when 7509 => DO <= x"00000000"; 
      when 7510 => DO <= x"00000000"; 
      when 7511 => DO <= x"00000000"; 
      when 7512 => DO <= x"00000000"; 
      when 7513 => DO <= x"00000000"; 
      when 7514 => DO <= x"00000000"; 
      when 7515 => DO <= x"00000000"; 
      when 7516 => DO <= x"00000000"; 
      when 7517 => DO <= x"00000000"; 
      when 7518 => DO <= x"00000000"; 
      when 7519 => DO <= x"00000000"; 
      when 7520 => DO <= x"00000000"; 
      when 7521 => DO <= x"00000000"; 
      when 7522 => DO <= x"00000000"; 
      when 7523 => DO <= x"00000000"; 
      when 7524 => DO <= x"00000000"; 
      when 7525 => DO <= x"00000000"; 
      when 7526 => DO <= x"00000000"; 
      when 7527 => DO <= x"00000000"; 
      when 7528 => DO <= x"00000000"; 
      when 7529 => DO <= x"00000000"; 
      when 7530 => DO <= x"00000000"; 
      when 7531 => DO <= x"00000000"; 
      when 7532 => DO <= x"00000000"; 
      when 7533 => DO <= x"00000000"; 
      when 7534 => DO <= x"00000000"; 
      when 7535 => DO <= x"00000000"; 
      when 7536 => DO <= x"00000000"; 
      when 7537 => DO <= x"00000000"; 
      when 7538 => DO <= x"00000000"; 
      when 7539 => DO <= x"00000000"; 
      when 7540 => DO <= x"00000000"; 
      when 7541 => DO <= x"00000000"; 
      when 7542 => DO <= x"00000000"; 
      when 7543 => DO <= x"00000000"; 
      when 7544 => DO <= x"00000000"; 
      when 7545 => DO <= x"00000000"; 
      when 7546 => DO <= x"00000000"; 
      when 7547 => DO <= x"00000000"; 
      when 7548 => DO <= x"00000000"; 
      when 7549 => DO <= x"00000000"; 
      when 7550 => DO <= x"00000000"; 
      when 7551 => DO <= x"00000000"; 
      when 7552 => DO <= x"00000000"; 
      when 7553 => DO <= x"00000000"; 
      when 7554 => DO <= x"00000000"; 
      when 7555 => DO <= x"00000000"; 
      when 7556 => DO <= x"00000000"; 
      when 7557 => DO <= x"00000000"; 
      when 7558 => DO <= x"00000000"; 
      when 7559 => DO <= x"00000000"; 
      when 7560 => DO <= x"00000000"; 
      when 7561 => DO <= x"00000000"; 
      when 7562 => DO <= x"00000000"; 
      when 7563 => DO <= x"00000000"; 
      when 7564 => DO <= x"00000000"; 
      when 7565 => DO <= x"00000000"; 
      when 7566 => DO <= x"00000000"; 
      when 7567 => DO <= x"00000000"; 
      when 7568 => DO <= x"00000000"; 
      when 7569 => DO <= x"00000000"; 
      when 7570 => DO <= x"00000000"; 
      when 7571 => DO <= x"00000000"; 
      when 7572 => DO <= x"00000000"; 
      when 7573 => DO <= x"00000000"; 
      when 7574 => DO <= x"00000000"; 
      when 7575 => DO <= x"00000000"; 
      when 7576 => DO <= x"00000000"; 
      when 7577 => DO <= x"00000000"; 
      when 7578 => DO <= x"00000000"; 
      when 7579 => DO <= x"00000000"; 
      when 7580 => DO <= x"00000000"; 
      when 7581 => DO <= x"00000000"; 
      when 7582 => DO <= x"00000000"; 
      when 7583 => DO <= x"00000000"; 
      when 7584 => DO <= x"00000000"; 
      when 7585 => DO <= x"00000000"; 
      when 7586 => DO <= x"00000000"; 
      when 7587 => DO <= x"00000000"; 
      when 7588 => DO <= x"00000000"; 
      when 7589 => DO <= x"00000000"; 
      when 7590 => DO <= x"00000000"; 
      when 7591 => DO <= x"00000000"; 
      when 7592 => DO <= x"00000000"; 
      when 7593 => DO <= x"00000000"; 
      when 7594 => DO <= x"00000000"; 
      when 7595 => DO <= x"00000000"; 
      when 7596 => DO <= x"00000000"; 
      when 7597 => DO <= x"00000000"; 
      when 7598 => DO <= x"00000000"; 
      when 7599 => DO <= x"00000000"; 
      when 7600 => DO <= x"00000000"; 
      when 7601 => DO <= x"00000000"; 
      when 7602 => DO <= x"00000000"; 
      when 7603 => DO <= x"00000000"; 
      when 7604 => DO <= x"00000000"; 
      when 7605 => DO <= x"00000000"; 
      when 7606 => DO <= x"00000000"; 
      when 7607 => DO <= x"00000000"; 
      when 7608 => DO <= x"00000000"; 
      when 7609 => DO <= x"00000000"; 
      when 7610 => DO <= x"00000000"; 
      when 7611 => DO <= x"00000000"; 
      when 7612 => DO <= x"00000000"; 
      when 7613 => DO <= x"00000000"; 
      when 7614 => DO <= x"00000000"; 
      when 7615 => DO <= x"00000000"; 
      when 7616 => DO <= x"00000000"; 
      when 7617 => DO <= x"00000000"; 
      when 7618 => DO <= x"00000000"; 
      when 7619 => DO <= x"00000000"; 
      when 7620 => DO <= x"00000000"; 
      when 7621 => DO <= x"00000000"; 
      when 7622 => DO <= x"00000000"; 
      when 7623 => DO <= x"00000000"; 
      when 7624 => DO <= x"00000000"; 
      when 7625 => DO <= x"00000000"; 
      when 7626 => DO <= x"00000000"; 
      when 7627 => DO <= x"00000000"; 
      when 7628 => DO <= x"00000000"; 
      when 7629 => DO <= x"00000000"; 
      when 7630 => DO <= x"00000000"; 
      when 7631 => DO <= x"00000000"; 
      when 7632 => DO <= x"00000000"; 
      when 7633 => DO <= x"00000000"; 
      when 7634 => DO <= x"00000000"; 
      when 7635 => DO <= x"00000000"; 
      when 7636 => DO <= x"00000000"; 
      when 7637 => DO <= x"00000000"; 
      when 7638 => DO <= x"00000000"; 
      when 7639 => DO <= x"00000000"; 
      when 7640 => DO <= x"00000000"; 
      when 7641 => DO <= x"00000000"; 
      when 7642 => DO <= x"00000000"; 
      when 7643 => DO <= x"00000000"; 
      when 7644 => DO <= x"00000000"; 
      when 7645 => DO <= x"00000000"; 
      when 7646 => DO <= x"00000000"; 
      when 7647 => DO <= x"00000000"; 
      when 7648 => DO <= x"00000000"; 
      when 7649 => DO <= x"00000000"; 
      when 7650 => DO <= x"00000000"; 
      when 7651 => DO <= x"00000000"; 
      when 7652 => DO <= x"00000000"; 
      when 7653 => DO <= x"00000000"; 
      when 7654 => DO <= x"00000000"; 
      when 7655 => DO <= x"00000000"; 
      when 7656 => DO <= x"00000000"; 
      when 7657 => DO <= x"00000000"; 
      when 7658 => DO <= x"00000000"; 
      when 7659 => DO <= x"00000000"; 
      when 7660 => DO <= x"00000000"; 
      when 7661 => DO <= x"00000000"; 
      when 7662 => DO <= x"00000000"; 
      when 7663 => DO <= x"00000000"; 
      when 7664 => DO <= x"00000000"; 
      when 7665 => DO <= x"00000000"; 
      when 7666 => DO <= x"00000000"; 
      when 7667 => DO <= x"00000000"; 
      when 7668 => DO <= x"00000000"; 
      when 7669 => DO <= x"00000000"; 
      when 7670 => DO <= x"00000000"; 
      when 7671 => DO <= x"00000000"; 
      when 7672 => DO <= x"00000000"; 
      when 7673 => DO <= x"00000000"; 
      when 7674 => DO <= x"00000000"; 
      when 7675 => DO <= x"00000000"; 
      when 7676 => DO <= x"00000000"; 
      when 7677 => DO <= x"00000000"; 
      when 7678 => DO <= x"00000000"; 
      when 7679 => DO <= x"00000000"; 
      when 7680 => DO <= x"00000000"; 
      when 7681 => DO <= x"00000000"; 
      when 7682 => DO <= x"00000000"; 
      when 7683 => DO <= x"00000000"; 
      when 7684 => DO <= x"00000000"; 
      when 7685 => DO <= x"00000000"; 
      when 7686 => DO <= x"00000000"; 
      when 7687 => DO <= x"00000000"; 
      when 7688 => DO <= x"00000000"; 
      when 7689 => DO <= x"00000000"; 
      when 7690 => DO <= x"00000000"; 
      when 7691 => DO <= x"00000000"; 
      when 7692 => DO <= x"00000000"; 
      when 7693 => DO <= x"00000000"; 
      when 7694 => DO <= x"00000000"; 
      when 7695 => DO <= x"00000000"; 
      when 7696 => DO <= x"00000000"; 
      when 7697 => DO <= x"00000000"; 
      when 7698 => DO <= x"00000000"; 
      when 7699 => DO <= x"00000000"; 
      when 7700 => DO <= x"00000000"; 
      when 7701 => DO <= x"00000000"; 
      when 7702 => DO <= x"00000000"; 
      when 7703 => DO <= x"00000000"; 
      when 7704 => DO <= x"00000000"; 
      when 7705 => DO <= x"00000000"; 
      when 7706 => DO <= x"00000000"; 
      when 7707 => DO <= x"00000000"; 
      when 7708 => DO <= x"00000000"; 
      when 7709 => DO <= x"00000000"; 
      when 7710 => DO <= x"00000000"; 
      when 7711 => DO <= x"00000000"; 
      when 7712 => DO <= x"00000000"; 
      when 7713 => DO <= x"00000000"; 
      when 7714 => DO <= x"00000000"; 
      when 7715 => DO <= x"00000000"; 
      when 7716 => DO <= x"00000000"; 
      when 7717 => DO <= x"00000000"; 
      when 7718 => DO <= x"00000000"; 
      when 7719 => DO <= x"00000000"; 
      when 7720 => DO <= x"00000000"; 
      when 7721 => DO <= x"00000000"; 
      when 7722 => DO <= x"00000000"; 
      when 7723 => DO <= x"00000000"; 
      when 7724 => DO <= x"00000000"; 
      when 7725 => DO <= x"00000000"; 
      when 7726 => DO <= x"00000000"; 
      when 7727 => DO <= x"00000000"; 
      when 7728 => DO <= x"00000000"; 
      when 7729 => DO <= x"00000000"; 
      when 7730 => DO <= x"00000000"; 
      when 7731 => DO <= x"00000000"; 
      when 7732 => DO <= x"00000000"; 
      when 7733 => DO <= x"00000000"; 
      when 7734 => DO <= x"00000000"; 
      when 7735 => DO <= x"00000000"; 
      when 7736 => DO <= x"00000000"; 
      when 7737 => DO <= x"00000000"; 
      when 7738 => DO <= x"00000000"; 
      when 7739 => DO <= x"00000000"; 
      when 7740 => DO <= x"00000000"; 
      when 7741 => DO <= x"00000000"; 
      when 7742 => DO <= x"00000000"; 
      when 7743 => DO <= x"00000000"; 
      when 7744 => DO <= x"00000000"; 
      when 7745 => DO <= x"00000000"; 
      when 7746 => DO <= x"00000000"; 
      when 7747 => DO <= x"00000000"; 
      when 7748 => DO <= x"00000000"; 
      when 7749 => DO <= x"00000000"; 
      when 7750 => DO <= x"00000000"; 
      when 7751 => DO <= x"00000000"; 
      when 7752 => DO <= x"00000000"; 
      when 7753 => DO <= x"00000000"; 
      when 7754 => DO <= x"00000000"; 
      when 7755 => DO <= x"00000000"; 
      when 7756 => DO <= x"00000000"; 
      when 7757 => DO <= x"00000000"; 
      when 7758 => DO <= x"00000000"; 
      when 7759 => DO <= x"00000000"; 
      when 7760 => DO <= x"00000000"; 
      when 7761 => DO <= x"00000000"; 
      when 7762 => DO <= x"00000000"; 
      when 7763 => DO <= x"00000000"; 
      when 7764 => DO <= x"00000000"; 
      when 7765 => DO <= x"00000000"; 
      when 7766 => DO <= x"00000000"; 
      when 7767 => DO <= x"00000000"; 
      when 7768 => DO <= x"00000000"; 
      when 7769 => DO <= x"00000000"; 
      when 7770 => DO <= x"00000000"; 
      when 7771 => DO <= x"00000000"; 
      when 7772 => DO <= x"00000000"; 
      when 7773 => DO <= x"00000000"; 
      when 7774 => DO <= x"00000000"; 
      when 7775 => DO <= x"00000000"; 
      when 7776 => DO <= x"00000000"; 
      when 7777 => DO <= x"00000000"; 
      when 7778 => DO <= x"00000000"; 
      when 7779 => DO <= x"00000000"; 
      when 7780 => DO <= x"00000000"; 
      when 7781 => DO <= x"00000000"; 
      when 7782 => DO <= x"00000000"; 
      when 7783 => DO <= x"00000000"; 
      when 7784 => DO <= x"00000000"; 
      when 7785 => DO <= x"00000000"; 
      when 7786 => DO <= x"00000000"; 
      when 7787 => DO <= x"00000000"; 
      when 7788 => DO <= x"00000000"; 
      when 7789 => DO <= x"00000000"; 
      when 7790 => DO <= x"00000000"; 
      when 7791 => DO <= x"00000000"; 
      when 7792 => DO <= x"00000000"; 
      when 7793 => DO <= x"00000000"; 
      when 7794 => DO <= x"00000000"; 
      when 7795 => DO <= x"00000000"; 
      when 7796 => DO <= x"00000000"; 
      when 7797 => DO <= x"00000000"; 
      when 7798 => DO <= x"00000000"; 
      when 7799 => DO <= x"00000000"; 
      when 7800 => DO <= x"00000000"; 
      when 7801 => DO <= x"00000000"; 
      when 7802 => DO <= x"00000000"; 
      when 7803 => DO <= x"00000000"; 
      when 7804 => DO <= x"00000000"; 
      when 7805 => DO <= x"00000000"; 
      when 7806 => DO <= x"00000000"; 
      when 7807 => DO <= x"00000000"; 
      when 7808 => DO <= x"00000000"; 
      when 7809 => DO <= x"00000000"; 
      when 7810 => DO <= x"00000000"; 
      when 7811 => DO <= x"00000000"; 
      when 7812 => DO <= x"00000000"; 
      when 7813 => DO <= x"00000000"; 
      when 7814 => DO <= x"00000000"; 
      when 7815 => DO <= x"00000000"; 
      when 7816 => DO <= x"00000000"; 
      when 7817 => DO <= x"00000000"; 
      when 7818 => DO <= x"00000000"; 
      when 7819 => DO <= x"00000000"; 
      when 7820 => DO <= x"00000000"; 
      when 7821 => DO <= x"00000000"; 
      when 7822 => DO <= x"00000000"; 
      when 7823 => DO <= x"00000000"; 
      when 7824 => DO <= x"00000000"; 
      when 7825 => DO <= x"00000000"; 
      when 7826 => DO <= x"00000000"; 
      when 7827 => DO <= x"00000000"; 
      when 7828 => DO <= x"00000000"; 
      when 7829 => DO <= x"00000000"; 
      when 7830 => DO <= x"00000000"; 
      when 7831 => DO <= x"00000000"; 
      when 7832 => DO <= x"00000000"; 
      when 7833 => DO <= x"00000000"; 
      when 7834 => DO <= x"00000000"; 
      when 7835 => DO <= x"00000000"; 
      when 7836 => DO <= x"00000000"; 
      when 7837 => DO <= x"00000000"; 
      when 7838 => DO <= x"00000000"; 
      when 7839 => DO <= x"00000000"; 
      when 7840 => DO <= x"00000000"; 
      when 7841 => DO <= x"00000000"; 
      when 7842 => DO <= x"00000000"; 
      when 7843 => DO <= x"00000000"; 
      when 7844 => DO <= x"00000000"; 
      when 7845 => DO <= x"00000000"; 
      when 7846 => DO <= x"00000000"; 
      when 7847 => DO <= x"00000000"; 
      when 7848 => DO <= x"00000000"; 
      when 7849 => DO <= x"00000000"; 
      when 7850 => DO <= x"00000000"; 
      when 7851 => DO <= x"00000000"; 
      when 7852 => DO <= x"00000000"; 
      when 7853 => DO <= x"00000000"; 
      when 7854 => DO <= x"00000000"; 
      when 7855 => DO <= x"00000000"; 
      when 7856 => DO <= x"00000000"; 
      when 7857 => DO <= x"00000000"; 
      when 7858 => DO <= x"00000000"; 
      when 7859 => DO <= x"00000000"; 
      when 7860 => DO <= x"00000000"; 
      when 7861 => DO <= x"00000000"; 
      when 7862 => DO <= x"00000000"; 
      when 7863 => DO <= x"00000000"; 
      when 7864 => DO <= x"00000000"; 
      when 7865 => DO <= x"00000000"; 
      when 7866 => DO <= x"00000000"; 
      when 7867 => DO <= x"00000000"; 
      when 7868 => DO <= x"00000000"; 
      when 7869 => DO <= x"00000000"; 
      when 7870 => DO <= x"00000000"; 
      when 7871 => DO <= x"00000000"; 
      when 7872 => DO <= x"00000000"; 
      when 7873 => DO <= x"00000000"; 
      when 7874 => DO <= x"00000000"; 
      when 7875 => DO <= x"00000000"; 
      when 7876 => DO <= x"00000000"; 
      when 7877 => DO <= x"00000000"; 
      when 7878 => DO <= x"00000000"; 
      when 7879 => DO <= x"00000000"; 
      when 7880 => DO <= x"00000000"; 
      when 7881 => DO <= x"00000000"; 
      when 7882 => DO <= x"00000000"; 
      when 7883 => DO <= x"00000000"; 
      when 7884 => DO <= x"00000000"; 
      when 7885 => DO <= x"00000000"; 
      when 7886 => DO <= x"00000000"; 
      when 7887 => DO <= x"00000000"; 
      when 7888 => DO <= x"00000000"; 
      when 7889 => DO <= x"00000000"; 
      when 7890 => DO <= x"00000000"; 
      when 7891 => DO <= x"00000000"; 
      when 7892 => DO <= x"00000000"; 
      when 7893 => DO <= x"00000000"; 
      when 7894 => DO <= x"00000000"; 
      when 7895 => DO <= x"00000000"; 
      when 7896 => DO <= x"00000000"; 
      when 7897 => DO <= x"00000000"; 
      when 7898 => DO <= x"00000000"; 
      when 7899 => DO <= x"00000000"; 
      when 7900 => DO <= x"00000000"; 
      when 7901 => DO <= x"00000000"; 
      when 7902 => DO <= x"00000000"; 
      when 7903 => DO <= x"00000000"; 
      when 7904 => DO <= x"00000000"; 
      when 7905 => DO <= x"00000000"; 
      when 7906 => DO <= x"00000000"; 
      when 7907 => DO <= x"00000000"; 
      when 7908 => DO <= x"00000000"; 
      when 7909 => DO <= x"00000000"; 
      when 7910 => DO <= x"00000000"; 
      when 7911 => DO <= x"00000000"; 
      when 7912 => DO <= x"00000000"; 
      when 7913 => DO <= x"00000000"; 
      when 7914 => DO <= x"00000000"; 
      when 7915 => DO <= x"00000000"; 
      when 7916 => DO <= x"00000000"; 
      when 7917 => DO <= x"00000000"; 
      when 7918 => DO <= x"00000000"; 
      when 7919 => DO <= x"00000000"; 
      when 7920 => DO <= x"00000000"; 
      when 7921 => DO <= x"00000000"; 
      when 7922 => DO <= x"00000000"; 
      when 7923 => DO <= x"00000000"; 
      when 7924 => DO <= x"00000000"; 
      when 7925 => DO <= x"00000000"; 
      when 7926 => DO <= x"00000000"; 
      when 7927 => DO <= x"00000000"; 
      when 7928 => DO <= x"00000000"; 
      when 7929 => DO <= x"00000000"; 
      when 7930 => DO <= x"00000000"; 
      when 7931 => DO <= x"00000000"; 
      when 7932 => DO <= x"00000000"; 
      when 7933 => DO <= x"00000000"; 
      when 7934 => DO <= x"00000000"; 
      when 7935 => DO <= x"00000000"; 
      when 7936 => DO <= x"00000000"; 
      when 7937 => DO <= x"00000000"; 
      when 7938 => DO <= x"00000000"; 
      when 7939 => DO <= x"00000000"; 
      when 7940 => DO <= x"00000000"; 
      when 7941 => DO <= x"00000000"; 
      when 7942 => DO <= x"00000000"; 
      when 7943 => DO <= x"00000000"; 
      when 7944 => DO <= x"00000000"; 
      when 7945 => DO <= x"00000000"; 
      when 7946 => DO <= x"00000000"; 
      when 7947 => DO <= x"00000000"; 
      when 7948 => DO <= x"00000000"; 
      when 7949 => DO <= x"00000000"; 
      when 7950 => DO <= x"00000000"; 
      when 7951 => DO <= x"00000000"; 
      when 7952 => DO <= x"00000000"; 
      when 7953 => DO <= x"00000000"; 
      when 7954 => DO <= x"00000000"; 
      when 7955 => DO <= x"00000000"; 
      when 7956 => DO <= x"00000000"; 
      when 7957 => DO <= x"00000000"; 
      when 7958 => DO <= x"00000000"; 
      when 7959 => DO <= x"00000000"; 
      when 7960 => DO <= x"00000000"; 
      when 7961 => DO <= x"00000000"; 
      when 7962 => DO <= x"00000000"; 
      when 7963 => DO <= x"00000000"; 
      when 7964 => DO <= x"00000000"; 
      when 7965 => DO <= x"00000000"; 
      when 7966 => DO <= x"00000000"; 
      when 7967 => DO <= x"00000000"; 
      when 7968 => DO <= x"00000000"; 
      when 7969 => DO <= x"00000000"; 
      when 7970 => DO <= x"00000000"; 
      when 7971 => DO <= x"00000000"; 
      when 7972 => DO <= x"00000000"; 
      when 7973 => DO <= x"00000000"; 
      when 7974 => DO <= x"00000000"; 
      when 7975 => DO <= x"00000000"; 
      when 7976 => DO <= x"00000000"; 
      when 7977 => DO <= x"00000000"; 
      when 7978 => DO <= x"00000000"; 
      when 7979 => DO <= x"00000000"; 
      when 7980 => DO <= x"00000000"; 
      when 7981 => DO <= x"00000000"; 
      when 7982 => DO <= x"00000000"; 
      when 7983 => DO <= x"00000000"; 
      when 7984 => DO <= x"00000000"; 
      when 7985 => DO <= x"00000000"; 
      when 7986 => DO <= x"00000000"; 
      when 7987 => DO <= x"00000000"; 
      when 7988 => DO <= x"00000000"; 
      when 7989 => DO <= x"00000000"; 
      when 7990 => DO <= x"00000000"; 
      when 7991 => DO <= x"00000000"; 
      when 7992 => DO <= x"00000000"; 
      when 7993 => DO <= x"00000000"; 
      when 7994 => DO <= x"00000000"; 
      when 7995 => DO <= x"00000000"; 
      when 7996 => DO <= x"00000000"; 
      when 7997 => DO <= x"00000000"; 
      when 7998 => DO <= x"00000000"; 
      when 7999 => DO <= x"00000000"; 
      when 8000 => DO <= x"00000000"; 
      when 8001 => DO <= x"00000000"; 
      when 8002 => DO <= x"00000000"; 
      when 8003 => DO <= x"00000000"; 
      when 8004 => DO <= x"00000000"; 
      when 8005 => DO <= x"00000000"; 
      when 8006 => DO <= x"00000000"; 
      when 8007 => DO <= x"00000000"; 
      when 8008 => DO <= x"00000000"; 
      when 8009 => DO <= x"00000000"; 
      when 8010 => DO <= x"00000000"; 
      when 8011 => DO <= x"00000000"; 
      when 8012 => DO <= x"00000000"; 
      when 8013 => DO <= x"00000000"; 
      when 8014 => DO <= x"00000000"; 
      when 8015 => DO <= x"00000000"; 
      when 8016 => DO <= x"00000000"; 
      when 8017 => DO <= x"00000000"; 
      when 8018 => DO <= x"00000000"; 
      when 8019 => DO <= x"00000000"; 
      when 8020 => DO <= x"00000000"; 
      when 8021 => DO <= x"00000000"; 
      when 8022 => DO <= x"00000000"; 
      when 8023 => DO <= x"00000000"; 
      when 8024 => DO <= x"00000000"; 
      when 8025 => DO <= x"00000000"; 
      when 8026 => DO <= x"00000000"; 
      when 8027 => DO <= x"00000000"; 
      when 8028 => DO <= x"00000000"; 
      when 8029 => DO <= x"00000000"; 
      when 8030 => DO <= x"00000000"; 
      when 8031 => DO <= x"00000000"; 
      when 8032 => DO <= x"00000000"; 
      when 8033 => DO <= x"00000000"; 
      when 8034 => DO <= x"00000000"; 
      when 8035 => DO <= x"00000000"; 
      when 8036 => DO <= x"00000000"; 
      when 8037 => DO <= x"00000000"; 
      when 8038 => DO <= x"00000000"; 
      when 8039 => DO <= x"00000000"; 
      when 8040 => DO <= x"00000000"; 
      when 8041 => DO <= x"00000000"; 
      when 8042 => DO <= x"00000000"; 
      when 8043 => DO <= x"00000000"; 
      when 8044 => DO <= x"00000000"; 
      when 8045 => DO <= x"00000000"; 
      when 8046 => DO <= x"00000000"; 
      when 8047 => DO <= x"00000000"; 
      when 8048 => DO <= x"00000000"; 
      when 8049 => DO <= x"00000000"; 
      when 8050 => DO <= x"00000000"; 
      when 8051 => DO <= x"00000000"; 
      when 8052 => DO <= x"00000000"; 
      when 8053 => DO <= x"00000000"; 
      when 8054 => DO <= x"00000000"; 
      when 8055 => DO <= x"00000000"; 
      when 8056 => DO <= x"00000000"; 
      when 8057 => DO <= x"00000000"; 
      when 8058 => DO <= x"00000000"; 
      when 8059 => DO <= x"00000000"; 
      when 8060 => DO <= x"00000000"; 
      when 8061 => DO <= x"00000000"; 
      when 8062 => DO <= x"00000000"; 
      when 8063 => DO <= x"00000000"; 
      when 8064 => DO <= x"00000000"; 
      when 8065 => DO <= x"00000000"; 
      when 8066 => DO <= x"00000000"; 
      when 8067 => DO <= x"00000000"; 
      when 8068 => DO <= x"00000000"; 
      when 8069 => DO <= x"00000000"; 
      when 8070 => DO <= x"00000000"; 
      when 8071 => DO <= x"00000000"; 
      when 8072 => DO <= x"00000000"; 
      when 8073 => DO <= x"00000000"; 
      when 8074 => DO <= x"00000000"; 
      when 8075 => DO <= x"00000000"; 
      when 8076 => DO <= x"00000000"; 
      when 8077 => DO <= x"00000000"; 
      when 8078 => DO <= x"00000000"; 
      when 8079 => DO <= x"00000000"; 
      when 8080 => DO <= x"00000000"; 
      when 8081 => DO <= x"00000000"; 
      when 8082 => DO <= x"00000000"; 
      when 8083 => DO <= x"00000000"; 
      when 8084 => DO <= x"00000000"; 
      when 8085 => DO <= x"00000000"; 
      when 8086 => DO <= x"00000000"; 
      when 8087 => DO <= x"00000000"; 
      when 8088 => DO <= x"00000000"; 
      when 8089 => DO <= x"00000000"; 
      when 8090 => DO <= x"00000000"; 
      when 8091 => DO <= x"00000000"; 
      when 8092 => DO <= x"00000000"; 
      when 8093 => DO <= x"00000000"; 
      when 8094 => DO <= x"00000000"; 
      when 8095 => DO <= x"00000000"; 
      when 8096 => DO <= x"00000000"; 
      when 8097 => DO <= x"00000000"; 
      when 8098 => DO <= x"00000000"; 
      when 8099 => DO <= x"00000000"; 
      when 8100 => DO <= x"00000000"; 
      when 8101 => DO <= x"00000000"; 
      when 8102 => DO <= x"00000000"; 
      when 8103 => DO <= x"00000000"; 
      when 8104 => DO <= x"00000000"; 
      when 8105 => DO <= x"00000000"; 
      when 8106 => DO <= x"00000000"; 
      when 8107 => DO <= x"00000000"; 
      when 8108 => DO <= x"00000000"; 
      when 8109 => DO <= x"00000000"; 
      when 8110 => DO <= x"00000000"; 
      when 8111 => DO <= x"00000000"; 
      when 8112 => DO <= x"00000000"; 
      when 8113 => DO <= x"00000000"; 
      when 8114 => DO <= x"00000000"; 
      when 8115 => DO <= x"00000000"; 
      when 8116 => DO <= x"00000000"; 
      when 8117 => DO <= x"00000000"; 
      when 8118 => DO <= x"00000000"; 
      when 8119 => DO <= x"00000000"; 
      when 8120 => DO <= x"00000000"; 
      when 8121 => DO <= x"00000000"; 
      when 8122 => DO <= x"00000000"; 
      when 8123 => DO <= x"00000000"; 
      when 8124 => DO <= x"00000000"; 
      when 8125 => DO <= x"00000000"; 
      when 8126 => DO <= x"00000000"; 
      when 8127 => DO <= x"00000000"; 
      when 8128 => DO <= x"00000000"; 
      when 8129 => DO <= x"00000000"; 
      when 8130 => DO <= x"00000000"; 
      when 8131 => DO <= x"00000000"; 
      when 8132 => DO <= x"00000000"; 
      when 8133 => DO <= x"00000000"; 
      when 8134 => DO <= x"00000000"; 
      when 8135 => DO <= x"00000000"; 
      when 8136 => DO <= x"00000000"; 
      when 8137 => DO <= x"00000000"; 
      when 8138 => DO <= x"00000000"; 
      when 8139 => DO <= x"00000000"; 
      when 8140 => DO <= x"00000000"; 
      when 8141 => DO <= x"00000000"; 
      when 8142 => DO <= x"00000000"; 
      when 8143 => DO <= x"00000000"; 
      when 8144 => DO <= x"00000000"; 
      when 8145 => DO <= x"00000000"; 
      when 8146 => DO <= x"00000000"; 
      when 8147 => DO <= x"00000000"; 
      when 8148 => DO <= x"00000000"; 
      when 8149 => DO <= x"00000000"; 
      when 8150 => DO <= x"00000000"; 
      when 8151 => DO <= x"00000000"; 
      when 8152 => DO <= x"00000000"; 
      when 8153 => DO <= x"00000000"; 
      when 8154 => DO <= x"00000000"; 
      when 8155 => DO <= x"00000000"; 
      when 8156 => DO <= x"00000000"; 
      when 8157 => DO <= x"00000000"; 
      when 8158 => DO <= x"00000000"; 
      when 8159 => DO <= x"00000000"; 
      when 8160 => DO <= x"00000000"; 
      when 8161 => DO <= x"00000000"; 
      when 8162 => DO <= x"00000000"; 
      when 8163 => DO <= x"00000000"; 
      when 8164 => DO <= x"00000000"; 
      when 8165 => DO <= x"00000000"; 
      when 8166 => DO <= x"00000000"; 
      when 8167 => DO <= x"00000000"; 
      when 8168 => DO <= x"00000000"; 
      when 8169 => DO <= x"00000000"; 
      when 8170 => DO <= x"00000000"; 
      when 8171 => DO <= x"00000000"; 
      when 8172 => DO <= x"00000000"; 
      when 8173 => DO <= x"00000000"; 
      when 8174 => DO <= x"00000000"; 
      when 8175 => DO <= x"00000000"; 
      when 8176 => DO <= x"00000000"; 
      when 8177 => DO <= x"00000000"; 
      when 8178 => DO <= x"00000000"; 
      when 8179 => DO <= x"00000000"; 
      when 8180 => DO <= x"00000000"; 
      when 8181 => DO <= x"00000000"; 
      when 8182 => DO <= x"00000000"; 
      when 8183 => DO <= x"00000000"; 
      when 8184 => DO <= x"00000000"; 
      when 8185 => DO <= x"00000000"; 
      when 8186 => DO <= x"00000000"; 
      when 8187 => DO <= x"00000000"; 
      when 8188 => DO <= x"00000000"; 
      when 8189 => DO <= x"00000000"; 
      when 8190 => DO <= x"00000000"; 
      when 8191 => DO <= x"00000000"; 
when others =>
end case;
end if;
end if;
end process;
end behave;
