library IEEE;
use IEEE.std_logic_1164.all; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.all;

entity internalram is
  port (
    CLKA:              in std_logic;
    WEA:  in std_logic;
    ENA:  in std_logic;
    MASKA:    in std_logic_vector(3 downto 0);
    ADDRA:         in std_logic_vector(14 downto 2);
    DIA:        in std_logic_vector(31 downto 0);
    DOA:         out std_logic_vector(31 downto 0);
    CLKB:              in std_logic;
    WEB:  in std_logic;
    ENB:  in std_logic;
    ADDRB:         in std_logic_vector(14 downto 2);
    DIB:        in std_logic_vector(31 downto 0);
    MASKB:    in std_logic_vector(3 downto 0);
    DOB:         out std_logic_vector(31 downto 0)
  );
end entity internalram;

architecture behave of internalram is

  subtype RAM_WORD is STD_LOGIC_VECTOR (7 downto 0);
  type RAM_TABLE is array (0 to 8191) of RAM_WORD;
 shared variable RAM0: RAM_TABLE := RAM_TABLE'(
x"00",x"61",x"bd",x"0a",x"a4",x"04",x"01",x"21",x"00",x"31",x"81",x"3f",x"10",x"63",x"02",x"00",x"03",x"52",x"14",x"42",x"ff",x"00",x"00",x"00",x"2d",x"21",x"10",x"02",x"60",x"41",x"41",x"d0",x"e0",x"e0",x"00",x"df",x"14",x"10",x"0c",x"1c",x"11",x"01",x"31",x"c0",x"10",x"31",x"00",x"31",x"f2",x"12",x"12",x"31",x"60",x"10",x"10",x"18",x"76",x"16",x"86",x"36",x"38",x"08",x"40",x"10",x"33",x"72",x"04",x"1a",x"14",x"3e",x"38",x"c0",x"10",x"3e",x"10",x"60",x"10",x"10",x"18",x"28",x"38",x"12",x"14",x"3c",x"38",x"40",x"10",x"3c",x"10",x"38",x"18",x"25",x"00",x"41",x"21",x"15",x"00",x"03",x"2f",x"12",x"41",x"32",x"1c",x"6f",x"5f",x"4f",x"df",x"d0",x"00",x"df",x"0c",x"5f",x"25",x"04",x"ed",x"10",x"51",x"2d",x"10",x"01",x"04",x"08",x"0c",x"0f",x"10",x"e0",x"10",x"37",x"00",x"37",x"79",x"f7",x"79",x"81",x"88",x"88",x"87",x"32",x"02",x"02",x"22",x"01",x"10",x"31",x"02",x"02",x"10",x"df",x"0c",x"08",x"04",x"18",x"24",x"04",x"01",x"1f",x"80",x"10",x"01",x"ff",x"81",x"ff",x"fb",x"f3",x"07",x"1f",x"01",x"10",x"2f",x"54",x"f2",x"00",x"a0",x"94",x"b6",x"99",x"29",x"00",x"c0",x"44",x"04",x"00",x"a0",x"3a",x"54",x"04",x"01",x"60",x"10",x"10",x"09",x"20",x"10",x"10",x"40",x"49",x"05",x"00",x"54",x"24",x"05",x"ff",x"25",x"c0",x"10",x"17",x"04",x"9f",x"e2",x"9f",x"e0",x"29",x"22",x"e2",x"04",x"00",x"4f",x"22",x"e2",x"42",x"10",x"11",x"c0",x"10",x"49",x"92",x"80",x"02",x"62",x"0f",x"26",x"82",x"ff",x"3f",x"f2",x"32",x"14",x"1c",x"10",x"01",x"26",x"14",x"02",x"71",x"40",x"10",x"18",x"42",x"2d",x"10",x"1f",x"14",x"71",x"04",x"10",x"04",x"04",x"04",x"22",x"61",x"f1",x"00",x"20",x"05",x"00",x"ff",x"f1",x"56",x"04",x"02",x"20",x"10",x"06",x"ff",x"a0",x"2f",x"05",x"00",x"56",x"04",x"01",x"60",x"10",x"06",x"ff",x"65",x"60",x"10",x"00",x"14",x"15",x"11",x"ed",x"10",x"14",x"e0",x"10",x"10",x"27",x"31",x"37",x"21",x"03",x"27",x"51",x"01",x"00",x"15",x"06",x"00",x"ff",x"f1",x"02",x"04",x"11",x"1e",x"66",x"06",x"ff",x"ff",x"f1",x"04",x"08",x"4f",x"df",x"d0",x"13",x"02",x"01",x"60",x"10",x"10",x"60",x"10",x"00",x"72",x"04",x"02",x"60",x"10",x"10",x"03",x"ff",x"c0",x"03",x"00",x"22",x"73",x"77",x"27",x"00",x"60",x"33",x"40",x"10",x"10",x"d0",x"31",x"10",x"01",x"00",x"80",x"12",x"32",x"01",x"ff",x"21",x"10",x"21",x"10",x"19",x"df",x"0c",x"08",x"04",x"18",x"1c",x"20",x"80",x"10",x"01",x"01",x"03",x"9b",x"11",x"24",x"7f",x"8f",x"08",x"14",x"78",x"00",x"00",x"10",x"1b",x"14",x"80",x"10",x"e0",x"10",x"60",x"10",x"00",x"10",x"f8",x"92",x"a0",x"08",x"00",x"0b",x"00",x"29",x"b1",x"7f",x"07",x"00",x"c0",x"37",x"10",x"24",x"a0",x"10",x"b9",x"2f",x"1f",x"01",x"20",x"10",x"10",x"10",x"95",x"2b",x"19",x"3f",x"7f",x"7d",x"01",x"00",x"af",x"25",x"53",x"fa",x"10",x"af",x"68",x"43",x"80",x"10",x"28",x"ff",x"3f",x"1f",x"b9",x"bb",x"0b",x"00",x"60",x"7f",x"72",x"ff",x"3f",x"80",x"3f",x"0b",x"14",x"8f",x"20",x"10",x"14",x"01",x"20",x"01",x"20",x"28",x"a0",x"10",x"04",x"08",x"0c",x"cf",x"10",x"f8",x"21",x"04",x"04",x"04",x"04",x"33",x"21",x"d0",x"31",x"72",x"71",x"32",x"32",x"12",x"10",x"8f",x"4f",x"24",x"5f",x"6f",x"3f",x"ed",x"10",x"fe",x"04",x"08",x"92",x"24",x"17",x"14",x"31",x"80",x"03",x"93",x"31",x"40",x"10",x"04",x"10",x"00",x"10",x"4e",x"0a",x"08",x"f8",x"74",x"87",x"ff",x"f8",x"b7",x"14",x"09",x"c0",x"09",x"10",x"00",x"3f",x"ff",x"f9",x"39",x"08",x"80",x"10",x"04",x"c0",x"10",x"75",x"5a",x"a9",x"55",x"53",x"05",x"08",x"06",x"25",x"f3",x"84",x"04",x"67",x"02",x"2f",x"1a",x"20",x"10",x"26",x"40",x"10",x"14",x"10",x"00",x"23",x"52",x"53",x"17",x"07",x"3f",x"01",x"e0",x"10",x"08",x"29",x"97",x"04",x"02",x"76",x"87",x"ff",x"41",x"01",x"6d",x"10",x"04",x"08",x"0c",x"8f",x"10",x"4f",x"af",x"07",x"89",x"a9",x"00",x"b4",x"10",x"ab",x"00",x"93",x"31",x"81",x"18",x"14",x"14",x"04",x"31",x"02",x"02",x"04",x"8f",x"10",x"df",x"0c",x"5f",x"6f",x"06",x"1c",x"3e",x"3c",x"3a",x"38",x"80",x"10",x"12",x"f8",x"24",x"6d",x"10",x"38",x"f2",x"f8",x"24",x"ed",x"10",x"38",x"60",x"10",x"3a",x"56",x"ff",x"6f",x"5f",x"4f",x"df",x"0f",x"10",x"4f",x"df",x"24",x"20",x"1c",x"28",x"30",x"f2",x"08",x"1f",x"21",x"00",x"68",x"33",x"11",x"16",x"1f",x"21",x"16",x"1f",x"31",x"16",x"1f",x"41",x"16",x"1f",x"51",x"16",x"73",x"40",x"10",x"3f",x"6f",x"16",x"00",x"80",x"1f",x"16",x"00",x"10",x"34",x"02",x"00",x"51",x"62",x"34",x"30",x"32",x"34",x"10",x"c0",x"10",x"32",x"01",x"00",x"1f",x"01",x"00",x"06",x"6f",x"6f",x"1f",x"1f",x"f2",x"04",x"00",x"54",x"38",x"30",x"32",x"42",x"05",x"32",x"08",x"1f",x"11",x"4f",x"3f",x"08",x"2f",x"22",x"08",x"3f",x"51",x"ff",x"f2",x"01",x"ed",x"10",x"00",x"54",x"1f",x"08",x"00",x"14",x"3c",x"00",x"50",x"20",x"10",x"42",x"14",x"32",x"40",x"00",x"44",x"00",x"4c",x"40",x"10",x"00",x"42",x"02",x"2f",x"08",x"00",x"2f",x"63",x"fb",x"1f",x"7f",x"21",x"01",x"00",x"1f",x"2f",x"11",x"22",x"03",x"00",x"48",x"40",x"28",x"48",x"0e",x"7f",x"41",x"01",x"00",x"1f",x"3f",x"12",x"48",x"13",x"1f",x"01",x"00",x"11",x"4c",x"c0",x"1f",x"a2",x"01",x"4c",x"31",x"f1",x"ed",x"10",x"31",x"ed",x"10",x"31",x"c6",x"7f",x"04",x"00",x"44",x"6d",x"10",x"01",x"00",x"05",x"00",x"44",x"00",x"03",x"2d",x"10",x"11",x"00",x"01",x"12",x"01",x"00",x"40",x"10",x"00",x"44",x"ed",x"10",x"01",x"00",x"12",x"6d",x"10",x"4c",x"21",x"1f",x"ad",x"10",x"30",x"00",x"4c",x"fc",x"6d",x"10",x"30",x"14",x"30",x"11",x"15",x"12",x"32",x"ad",x"10",x"1f",x"11",x"15",x"12",x"4a",x"ed",x"10",x"ff",x"f3",x"45",x"00",x"10",x"18",x"00",x"c0",x"91",x"0d",x"10",x"e0",x"55",x"c0",x"10",x"00",x"60",x"10",x"10",x"5e",x"15",x"32",x"10",x"4e",x"01",x"b1",x"cd",x"10",x"a0",x"f1",x"cd",x"10",x"a0",x"8a",x"25",x"01",x"21",x"0d",x"10",x"01",x"03",x"01",x"01",x"08",x"5f",x"08",x"4f",x"21",x"08",x"2f",x"02",x"06",x"12",x"00",x"50",x"5d",x"08",x"2f",x"42",x"21",x"08",x"1f",x"08",x"2f",x"08",x"3f",x"41",x"00",x"4c",x"01",x"05",x"15",x"11",x"20",x"01",x"00",x"01",x"10",x"3a",x"00",x"50",x"01",x"c0",x"10",x"5f",x"0d",x"10",x"40",x"15",x"25",x"23",x"03",x"00",x"35",x"08",x"7f",x"47",x"c0",x"10",x"5f",x"4d",x"10",x"40",x"15",x"25",x"43",x"02",x"00",x"35",x"08",x"2f",x"42",x"80",x"10",x"5f",x"8d",x"10",x"40",x"15",x"08",x"3f",x"08",x"2f",x"13",x"ff",x"f1",x"06",x"63",x"16",x"fe",x"08",x"4f",x"08",x"2f",x"08",x"5f",x"08",x"3f",x"08",x"5f",x"08",x"2f",x"08",x"4f",x"cd",x"10",x"00",x"48",x"5f",x"48",x"13",x"d1",x"42",x"13",x"41",x"2d",x"12",x"60",x"cd",x"10",x"ad",x"10",x"03",x"16",x"00",x"50",x"38",x"15",x"40",x"10",x"08",x"2f",x"61",x"04",x"36",x"11",x"40",x"10",x"51",x"00",x"5c",x"21",x"e0",x"10",x"63",x"4c",x"21",x"2d",x"10",x"51",x"2d",x"10",x"41",x"c4",x"3c",x"12",x"60",x"0d",x"10",x"ed",x"10",x"00",x"03",x"16",x"00",x"50",x"37",x"15",x"40",x"10",x"08",x"2f",x"61",x"80",x"04",x"36",x"f1",x"40",x"10",x"08",x"2f",x"08",x"3f",x"08",x"4f",x"51",x"06",x"21",x"e0",x"10",x"60",x"12",x"16",x"63",x"4c",x"21",x"11",x"0d",x"10",x"60",x"60",x"12",x"61",x"02",x"4d",x"10",x"60",x"61",x"11",x"a1",x"42",x"11",x"1f",x"12",x"02",x"00",x"08",x"6f",x"80",x"08",x"6f",x"25",x"60",x"10",x"00",x"4c",x"05",x"06",x"21",x"41",x"3a",x"61",x"11",x"16",x"00",x"16",x"15",x"60",x"10",x"50",x"63",x"12",x"c0",x"10",x"02",x"00",x"08",x"4f",x"02",x"63",x"41",x"01",x"31",x"11",x"cd",x"10",x"ff",x"f1",x"02",x"12",x"ff",x"1f",x"42",x"01",x"02",x"08",x"7f",x"20",x"10",x"a0",x"10",x"04",x"05",x"76",x"01",x"31",x"d1",x"0d",x"10",x"ff",x"f1",x"15",x"14",x"20",x"10",x"a0",x"10",x"06",x"05",x"74",x"01",x"31",x"91",x"0d",x"10",x"ff",x"f1",x"15",x"16",x"20",x"10",x"00",x"44",x"00",x"21",x"60",x"10",x"10",x"11",x"00",x"f1",x"40",x"10",x"61",x"10",x"08",x"1f",x"31",x"00",x"01",x"2f",x"11",x"01",x"41",x"14",x"00",x"5c",x"ed",x"10",x"41",x"c4",x"39",x"12",x"60",x"04",x"1f",x"f1",x"0d",x"10",x"61",x"61",x"0f",x"f1",x"60",x"01",x"0d",x"10",x"00",x"68",x"2a",x"6f",x"5f",x"4f",x"df",x"cf",x"d0",x"00",x"df",x"0c",x"08",x"71",x"41",x"31",x"11",x"04",x"ad",x"52",x"0f",x"5f",x"4f",x"df",x"d0",x"cf",x"28",x"4f",x"5f",x"15",x"6f",x"05",x"03",x"01",x"91",x"10",x"15",x"0a",x"07",x"5a",x"01",x"87",x"87",x"ff",x"11",x"80",x"10",x"15",x"0a",x"08",x"5a",x"02",x"01",x"e7",x"88",x"08",x"e0",x"10",x"51",x"ff",x"3f",x"01",x"0a",x"15",x"08",x"09",x"02",x"99",x"10",x"b3",x"00",x"a2",x"00",x"1b",x"40",x"10",x"b2",x"9a",x"60",x"10",x"9a",x"40",x"10",x"02",x"ad",x"10",x"14",x"06",x"61",x"65",x"03",x"e1",x"78",x"89",x"18",x"aa",x"49",x"99",x"99",x"9a",x"93",x"ff",x"16",x"56",x"ff",x"01",x"0b",x"15",x"09",x"0a",x"02",x"aa",x"10",x"67",x"00",x"a3",x"40",x"e6",x"ba",x"00",x"0e",x"6e",x"ab",x"20",x"10",x"ab",x"00",x"10",x"e6",x"0d",x"12",x"20",x"10",x"1c",x"6e",x"14",x"03",x"37",x"e6",x"0a",x"02",x"08",x"0e",x"0b",x"5a",x"bb",x"ee",x"2b",x"bb",x"bb",x"eb",x"b9",x"ff",x"17",x"98",x"40",x"10",x"51",x"ff",x"2f",x"01",x"0b",x"15",x"09",x"0a",x"02",x"aa",x"27",x"00",x"a3",x"40",x"e6",x"ba",x"00",x"0e",x"6e",x"ab",x"60",x"10",x"ab",x"40",x"10",x"1c",x"e6",x"0c",x"12",x"c0",x"10",x"2f",x"01",x"f7",x"18",x"14",x"08",x"1f",x"89",x"0b",x"02",x"0a",x"0a",x"01",x"01",x"11",x"e5",x"1e",x"91",x"01",x"11",x"12",x"21",x"22",x"31",x"21",x"1b",x"ff",x"ba",x"ef",x"59",x"ff",x"1f",x"11",x"a0",x"10",x"04",x"03",x"07",x"78",x"22",x"e2",x"2f",x"93",x"a0",x"10",x"03",x"10",x"a9",x"00",x"0b",x"18",x"58",x"ff",x"11",x"51",x"ff",x"2f",x"80",x"01",x"3f",x"ad",x"10",x"01",x"0b",x"12",x"04",x"0b",x"12",x"ad",x"10",x"40",x"10",x"28",x"14",x"25",x"07",x"08",x"57",x"01",x"98",x"09",x"60",x"10",x"52",x"ff",x"a0",x"01",x"0b",x"6f",x"5f",x"4f",x"df",x"4f",x"10",x"e0",x"10",x"71",x"09",x"0a",x"19",x"01",x"ba",x"ba",x"ff",x"17",x"80",x"10",x"10",x"cf",x"01",x"00",x"07",x"08",x"89",x"19",x"ba",x"bb",x"3b",x"bb",x"b4",x"ba",x"ff",x"17",x"e0",x"10",x"4f",x"10",x"07",x"04",x"01",x"00",x"08",x"04",x"81",x"0b",x"0e",x"02",x"ee",x"39",x"00",x"a7",x"00",x"15",x"40",x"10",x"57",x"e4",x"a0",x"10",x"e4",x"80",x"10",x"4f",x"71",x"d0",x"8f",x"04",x"01",x"00",x"07",x"02",x"0a",x"0b",x"08",x"05",x"01",x"1b",x"01",x"35",x"55",x"55",x"0e",x"a0",x"10",x"98",x"e0",x"10",x"4f",x"8f",x"10",x"4f",x"5f",x"6f",x"e0",x"10",x"71",x"09",x"0a",x"0e",x"02",x"0a",x"06",x"05",x"1e",x"55",x"66",x"35",x"55",x"55",x"65",x"5b",x"ff",x"19",x"19",x"ff",x"17",x"80",x"10",x"5f",x"4f",x"cf",x"10",x"4f",x"5f",x"6f",x"0c",x"00",x"10",x"f2",x"71",x"0b",x"10",x"0c",x"07",x"06",x"02",x"0e",x"61",x"a6",x"16",x"b8",x"01",x"01",x"48",x"88",x"88",x"07",x"05",x"02",x"97",x"07",x"40",x"10",x"5e",x"20",x"10",x"10",x"17",x"ff",x"6f",x"04",x"08",x"d0",x"00",x"17",x"4f",x"5f",x"6f",x"0c",x"40",x"10",x"f1",x"a0",x"10",x"31",x"01",x"09",x"03",x"c0",x"10",x"c3",x"32",x"03",x"00",x"17",x"91",x"05",x"86",x"00",x"0b",x"1f",x"10",x"ba",x"08",x"0a",x"15",x"0b",x"01",x"01",x"b2",x"68",x"b4",x"f4",x"16",x"4a",x"ff",x"19",x"19",x"ff",x"8f",x"37",x"33",x"27",x"04",x"78",x"28",x"18",x"5f",x"4f",x"0f",x"10",x"df",x"0c",x"08",x"6f",x"4f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"14",x"5f",x"15",x"60",x"10",x"10",x"50",x"30",x"01",x"11",x"f2",x"21",x"12",x"1f",x"11",x"60",x"10",x"10",x"60",x"5f",x"11",x"04",x"58",x"00",x"51",x"c2",x"00",x"62",x"31",x"a0",x"10",x"50",x"50",x"15",x"60",x"10",x"10",x"50",x"30",x"01",x"11",x"f2",x"21",x"12",x"1f",x"11",x"60",x"10",x"10",x"50",x"58",x"20",x"10",x"54",x"c1",x"00",x"21",x"65",x"a0",x"10",x"50",x"64",x"10",x"05",x"12",x"30",x"05",x"12",x"14",x"05",x"12",x"34",x"05",x"12",x"18",x"05",x"12",x"38",x"05",x"12",x"1c",x"05",x"12",x"3c",x"05",x"12",x"20",x"05",x"12",x"40",x"05",x"12",x"24",x"05",x"12",x"44",x"05",x"12",x"28",x"05",x"12",x"48",x"05",x"12",x"2c",x"05",x"12",x"4c",x"05",x"6f",x"5f",x"4f",x"df",x"d0",x"00",x"03",x"0a",x"00",x"40",x"10",x"f8",x"09",x"0b",x"80",x"10",x"01",x"33",x"00",x"03",x"00",x"23",x"00",x"60",x"10",x"d0",x"93",x"01",x"32",x"13",x"08",x"e0",x"10",x"a0",x"10",x"80",x"10",x"00",x"eb",x"01",x"32",x"13",x"10",x"e0",x"10",x"80",x"10",x"00",x"32",x"13",x"18",x"d0",x"0a",x"aa",x"01",x"a0",x"10",x"d0",x"0a",x"aa",x"00",x"23",x"c0",x"10",x"40",x"10",x"00",x"10",x"40",x"10",x"20",x"10",x"a0",x"10",x"20",x"10",x"0c",x"32",x"63",x"00",x"53",x"00",x"9a",x"83",x"20",x"10",x"14",x"32",x"33",x"10",x"20",x"10",x"d0",x"0a",x"aa",x"00",x"80",x"10",x"08",x"13",x"08",x"60",x"10",x"00",x"a3",x"83",x"43",x"e0",x"10",x"10",x"d0",x"0a",x"aa",x"00",x"e0",x"32",x"13",x"04",x"a2",x"a2",x"01",x"01",x"a0",x"10",x"13",x"fe",x"c0",x"7b",x"10",x"01",x"31",x"10",x"0c",x"32",x"80",x"32",x"13",x"04",x"10",x"10",x"32",x"c0",x"32",x"13",x"14",x"01",x"c0",x"cf",x"4f",x"5f",x"6f",x"1f",x"18",x"07",x"01",x"a0",x"1a",x"81",x"1a",x"04",x"05",x"01",x"80",x"10",x"00",x"06",x"20",x"10",x"0b",x"0a",x"16",x"aa",x"a0",x"10",x"53",x"9a",x"7a",x"a5",x"46",x"00",x"36",x"00",x"6a",x"2a",x"ff",x"40",x"6a",x"2a",x"00",x"76",x"ff",x"51",x"ca",x"0a",x"40",x"10",x"01",x"a1",x"5e",x"ff",x"51",x"ca",x"0a",x"1a",x"41",x"00",x"10",x"01",x"a1",x"5e",x"ff",x"1f",x"17",x"00",x"73",x"71",x"21",x"2d",x"10",x"04",x"08",x"0c",x"4f",x"10",x"01",x"60",x"10",x"60",x"10",x"10",x"63",x"10",x"60",x"10",x"60",x"10",x"10",x"63",x"10",x"00",x"10",x"63",x"10",x"63",x"10",x"80",x"10",x"63",x"d0",x"23",x"21",x"17",x"09",x"40",x"10",x"29",x"88",x"12",x"28",x"78",x"02",x"00",x"39",x"00",x"88",x"29",x"01",x"09",x"02",x"78",x"0a",x"00",x"39",x"88",x"9a",x"8a",x"18",x"a8",x"0a",x"40",x"10",x"29",x"0f",x"01",x"09",x"04",x"78",x"0a",x"00",x"39",x"88",x"9a",x"8a",x"18",x"a8",x"0a",x"40",x"10",x"29",x"0f",x"01",x"09",x"06",x"78",x"0a",x"00",x"39",x"11",x"99",x"91",x"0a",x"0f",x"97",x"00",x"37",x"11",x"22",x"21",x"00",x"21",x"10",x"df",x"04",x"f1",x"41",x"fe",x"12",x"08",x"fe",x"4f",x"df",x"d0",x"4f",x"4f",x"5f",x"14",x"00",x"01",x"fe",x"12",x"00",x"41",x"08",x"fe",x"12",x"10",x"8d",x"10",x"41",x"cd",x"10",x"04",x"08",x"cf",x"10",x"df",x"04",x"f1",x"41",x"fe",x"12",x"00",x"41",x"08",x"fe",x"4f",x"df",x"d0",x"01",x"10",x"71",x"37",x"40",x"10",x"d0",x"42",x"23",x"72",x"37",x"40",x"10",x"d0",x"4f",x"df",x"14",x"10",x"0c",x"00",x"2c",x"00",x"28",x"00",x"24",x"00",x"dc",x"f5",x"00",x"dc",x"00",x"d8",x"00",x"02",x"2f",x"12",x"00",x"04",x"10",x"01",x"52",x"08",x"0b",x"f9",x"aa",x"60",x"1b",x"31",x"12",x"33",x"60",x"10",x"60",x"10",x"10",x"21",x"10",x"40",x"10",x"60",x"10",x"10",x"21",x"10",x"c0",x"10",x"e0",x"41",x"10",x"80",x"10",x"a0",x"37",x"08",x"97",x"00",x"12",x"8a",x"33",x"83",x"d0",x"d0",x"97",x"00",x"10",x"10",x"93",x"40",x"10",x"00",x"d8",x"32",x"23",x"00",x"3f",x"82",x"02",x"c0",x"10",x"1b",x"81",x"32",x"e3",x"00",x"40",x"01",x"bf",x"01",x"8f",x"2b",x"32",x"37",x"97",x"07",x"80",x"10",x"3b",x"7a",x"22",x"72",x"d0",x"d0",x"98",x"00",x"10",x"10",x"00",x"f4",x"00",x"e8",x"00",x"e4",x"80",x"f7",x"08",x"60",x"10",x"00",x"d8",x"2b",x"33",x"37",x"00",x"7f",x"73",x"02",x"01",x"bf",x"07",x"00",x"76",x"32",x"c2",x"00",x"e0",x"01",x"1f",x"21",x"11",x"00",x"e4",x"40",x"32",x"a3",x"80",x"10",x"40",x"10",x"60",x"10",x"80",x"10",x"00",x"01",x"2f",x"01",x"01",x"2f",x"20",x"27",x"00",x"97",x"00",x"f7",x"00",x"c0",x"10",x"00",x"37",x"04",x"47",x"00",x"e0",x"10",x"00",x"f4",x"12",x"00",x"f4",x"10",x"80",x"10",x"20",x"10",x"80",x"10",x"04",x"03",x"00",x"d8",x"31",x"12",x"00",x"2f",x"21",x"00",x"f4",x"08",x"04",x"01",x"4f",x"0d",x"10",x"01",x"6f",x"20",x"10",x"00",x"f4",x"23",x"00",x"f4",x"10",x"80",x"10",x"04",x"01",x"5f",x"c3",x"c1",x"00",x"d8",x"32",x"04",x"00",x"d8",x"22",x"00",x"f8",x"00",x"e0",x"10",x"00",x"f4",x"00",x"e4",x"a2",x"a1",x"60",x"10",x"63",x"00",x"f8",x"a9",x"81",x"11",x"23",x"33",x"1f",x"3f",x"9f",x"3b",x"37",x"83",x"23",x"7f",x"33",x"1c",x"1d",x"02",x"04",x"27",x"77",x"1e",x"3f",x"9f",x"3b",x"37",x"83",x"23",x"7f",x"33",x"22",x"23",x"04",x"04",x"27",x"77",x"24",x"3f",x"9f",x"3b",x"37",x"83",x"32",x"7f",x"22",x"28",x"01",x"5f",x"a2",x"80",x"10",x"04",x"01",x"4f",x"24",x"00",x"00",x"10",x"51",x"43",x"15",x"1f",x"45",x"60",x"10",x"80",x"10",x"00",x"f1",x"e2",x"01",x"21",x"00",x"f8",x"00",x"ec",x"41",x"00",x"10",x"18",x"71",x"00",x"44",x"00",x"f1",x"42",x"00",x"e0",x"05",x"6d",x"10",x"62",x"61",x"15",x"2d",x"10",x"14",x"33",x"61",x"11",x"01",x"6d",x"10",x"00",x"e0",x"27",x"10",x"60",x"10",x"10",x"18",x"01",x"7f",x"71",x"41",x"33",x"a6",x"a2",x"11",x"41",x"34",x"01",x"7f",x"14",x"60",x"a6",x"f2",x"f1",x"42",x"62",x"21",x"00",x"ec",x"01",x"43",x"fe",x"01",x"2f",x"01",x"01",x"00",x"80",x"10",x"00",x"e8",x"00",x"f0",x"ff",x"80",x"10",x"05",x"71",x"51",x"01",x"7f",x"43",x"14",x"01",x"7f",x"45",x"00",x"e8",x"05",x"07",x"01",x"00",x"1f",x"c2",x"21",x"04",x"00",x"d8",x"00",x"e8",x"f3",x"00",x"02",x"00",x"f4",x"23",x"3f",x"6f",x"a0",x"10",x"00",x"e8",x"03",x"0c",x"15",x"05",x"01",x"2f",x"01",x"01",x"00",x"e0",x"10",x"00",x"e8",x"00",x"e4",x"ff",x"80",x"10",x"02",x"51",x"43",x"13",x"00",x"1f",x"c2",x"21",x"04",x"00",x"d8",x"02",x"11",x"80",x"10",x"a0",x"10",x"00",x"d8",x"23",x"21",x"12",x"00",x"d8",x"01",x"1f",x"00",x"1f",x"12",x"00",x"2f",x"01",x"7f",x"02",x"72",x"80",x"10",x"01",x"e2",x"00",x"f0",x"a0",x"10",x"92",x"00",x"10",x"00",x"e4",x"00",x"00",x"1f",x"c2",x"21",x"04",x"00",x"d8",x"08",x"00",x"38",x"18",x"01",x"00",x"81",x"06",x"00",x"14",x"11",x"01",x"00",x"f6",x"06",x"ff",x"01",x"2f",x"01",x"06",x"01",x"02",x"01",x"1f",x"16",x"00",x"c0",x"10",x"02",x"03",x"01",x"3f",x"01",x"8f",x"6d",x"10",x"00",x"e0",x"81",x"01",x"1f",x"01",x"1f",x"15",x"01",x"51",x"15",x"00",x"e4",x"01",x"00",x"e0",x"21",x"11",x"f7",x"15",x"21",x"e0",x"10",x"00",x"10",x"15",x"a0",x"10",x"00",x"e4",x"00",x"e8",x"10",x"00",x"e8",x"01",x"01",x"5f",x"c0",x"10",x"00",x"1f",x"c2",x"ff",x"31",x"12",x"00",x"2f",x"11",x"51",x"00",x"10",x"61",x"e0",x"10",x"00",x"f0",x"04",x"00",x"f4",x"04",x"00",x"f8",x"01",x"2f",x"01",x"1f",x"6d",x"10",x"01",x"00",x"05",x"00",x"f8",x"03",x"21",x"00",x"f8",x"00",x"e0",x"00",x"ec",x"1a",x"f1",x"40",x"10",x"01",x"3f",x"02",x"32",x"00",x"08",x"21",x"00",x"e4",x"92",x"00",x"f4",x"00",x"10",x"00",x"e0",x"00",x"d3",x"00",x"01",x"2f",x"01",x"1f",x"f1",x"01",x"41",x"00",x"01",x"00",x"00",x"10",x"1c",x"11",x"13",x"01",x"00",x"e8",x"03",x"01",x"01",x"f1",x"00",x"e8",x"c0",x"10",x"52",x"26",x"11",x"00",x"73",x"11",x"72",x"12",x"c0",x"10",x"01",x"1f",x"12",x"00",x"10",x"01",x"04",x"01",x"f4",x"24",x"19",x"01",x"1a",x"02",x"1b",x"03",x"1c",x"04",x"1d",x"05",x"1e",x"06",x"1f",x"07",x"20",x"08",x"21",x"09",x"22",x"0a",x"23",x"0b",x"24",x"0c",x"25",x"0d",x"26",x"0e",x"27",x"0f",x"28",x"10",x"11",x"00",x"e0",x"43",x"02",x"05",x"15",x"01",x"f4",x"01",x"1f",x"01",x"f7",x"00",x"f3",x"13",x"61",x"32",x"c0",x"10",x"16",x"00",x"11",x"01",x"1f",x"12",x"c0",x"10",x"71",x"04",x"02",x"6d",x"10",x"01",x"1f",x"11",x"f4",x"01",x"1f",x"b3",x"62",x"40",x"10",x"02",x"1f",x"21",x"91",x"71",x"80",x"10",x"20",x"71",x"02",x"8f",x"02",x"9f",x"01",x"3f",x"51",x"00",x"26",x"00",x"01",x"2f",x"20",x"10",x"00",x"00",x"c0",x"10",x"38",x"30",x"08",x"34",x"04",x"00",x"e0",x"00",x"ec",x"00",x"f8",x"ed",x"10",x"30",x"d1",x"00",x"21",x"04",x"25",x"f1",x"01",x"2f",x"53",x"f4",x"1f",x"f1",x"1f",x"01",x"3f",x"01",x"1f",x"01",x"2f",x"6d",x"10",x"34",x"c0",x"10",x"00",x"40",x"d2",x"00",x"88",x"00",x"04",x"15",x"02",x"8f",x"60",x"10",x"10",x"26",x"32",x"60",x"26",x"05",x"00",x"01",x"2f",x"63",x"11",x"11",x"13",x"20",x"10",x"08",x"00",x"51",x"02",x"00",x"14",x"1f",x"01",x"00",x"01",x"1f",x"01",x"2f",x"03",x"4d",x"10",x"01",x"00",x"04",x"10",x"ff",x"51",x"f4",x"00",x"e0",x"00",x"01",x"1f",x"d2",x"04",x"21",x"10",x"00",x"fc",x"61",x"41",x"ed",x"10",x"00",x"14",x"a2",x"04",x"6d",x"10",x"ed",x"10",x"42",x"03",x"00",x"e0",x"41",x"21",x"a2",x"23",x"01",x"05",x"00",x"08",x"84",x"00",x"f4",x"00",x"10",x"01",x"2f",x"01",x"00",x"02",x"00",x"00",x"00",x"40",x"12",x"47",x"00",x"07",x"00",x"e7",x"00",x"20",x"03",x"57",x"00",x"57",x"ff",x"27",x"01",x"01",x"e0",x"10",x"87",x"60",x"10",x"03",x"e0",x"10",x"07",x"03",x"87",x"e0",x"10",x"10",x"01",x"32",x"02",x"80",x"10",x"00",x"10",x"88",x"f2",x"72",x"07",x"00",x"03",x"12",x"c0",x"10",x"03",x"ff",x"03",x"80",x"10",x"10",x"12",x"07",x"00",x"57",x"00",x"57",x"ff",x"27",x"98",x"87",x"09",x"ff",x"e9",x"00",x"87",x"27",x"00",x"31",x"00",x"71",x"12",x"71",x"02",x"0a",x"00",x"1f",x"01",x"8f",x"02",x"9f",x"88",x"f2",x"01",x"01",x"e0",x"10",x"01",x"01",x"e0",x"10",x"17",x"60",x"10",x"05",x"59",x"82",x"80",x"10",x"60",x"10",x"10",x"00",x"01",x"6f",x"92",x"04",x"61",x"2d",x"10",x"00",x"f4",x"f4",x"00",x"f0",x"10",x"01",x"2f",x"f1",x"21",x"60",x"10",x"00",x"f0",x"11",x"00",x"f0",x"81",x"00",x"10",x"60",x"10",x"10",x"00",x"08",x"00",x"f0",x"00",x"12",x"6d",x"10",x"f4",x"00",x"f0",x"10",x"01",x"6f",x"01",x"2f",x"01",x"00",x"10",x"00",x"f0",x"10",x"88",x"f3",x"11",x"33",x"60",x"10",x"10",x"00",x"f0",x"15",x"e0",x"10",x"02",x"2d",x"10",x"61",x"a0",x"10",x"06",x"38",x"30",x"1f",x"f1",x"1f",x"01",x"1f",x"01",x"2f",x"8d",x"10",x"34",x"c0",x"10",x"00",x"40",x"d2",x"00",x"88",x"00",x"04",x"03",x"00",x"60",x"01",x"14",x"00",x"40",x"10",x"02",x"14",x"41",x"ad",x"10",x"01",x"02",x"fc",x"7f",x"02",x"00",x"10",x"08",x"07",x"01",x"24",x"60",x"10",x"10",x"14",x"3f",x"37",x"32",x"ff",x"21",x"c0",x"10",x"13",x"14",x"01",x"02",x"fc",x"80",x"7f",x"12",x"72",x"00",x"e3",x"14",x"34",x"31",x"03",x"fb",x"60",x"14",x"fb",x"01",x"00",x"2f",x"02",x"00",x"dc",x"f8",x"63",x"93",x"04",x"0a",x"ff",x"22",x"29",x"01",x"01",x"02",x"ff",x"6f",x"5f",x"4f",x"df",x"02",x"10",x"cf",x"4f",x"5f",x"6f",x"18",x"02",x"7c",x"12",x"80",x"10",x"21",x"02",x"62",x"01",x"00",x"fa",x"01",x"fe",x"20",x"10",x"02",x"01",x"00",x"f9",x"00",x"60",x"41",x"01",x"00",x"f4",x"80",x"01",x"d2",x"09",x"10",x"1c",x"11",x"12",x"71",x"03",x"04",x"8f",x"17",x"08",x"70",x"00",x"80",x"83",x"00",x"40",x"f4",x"5c",x"10",x"5c",x"10",x"5c",x"40",x"10",x"35",x"04",x"4f",x"7f",x"09",x"21",x"6c",x"00",x"06",x"af",x"f1",x"42",x"61",x"54",x"ad",x"10",x"58",x"11",x"54",x"51",x"2d",x"10",x"16",x"80",x"10",x"10",x"16",x"1f",x"6f",x"45",x"78",x"40",x"10",x"6f",x"1f",x"2f",x"4f",x"61",x"11",x"01",x"00",x"13",x"00",x"60",x"41",x"36",x"05",x"64",x"40",x"f3",x"5c",x"00",x"01",x"00",x"24",x"1f",x"37",x"c0",x"10",x"60",x"10",x"10",x"14",x"01",x"24",x"10",x"80",x"10",x"14",x"2f",x"5f",x"01",x"01",x"00",x"17",x"00",x"00",x"2f",x"f1",x"73",x"12",x"2d",x"10",x"f7",x"10",x"1f",x"15",x"00",x"46",x"04",x"75",x"43",x"05",x"57",x"58",x"64",x"e0",x"10",x"42",x"f3",x"01",x"33",x"12",x"ff",x"54",x"60",x"10",x"10",x"02",x"75",x"04",x"54",x"40",x"41",x"04",x"08",x"0c",x"4f",x"10",x"17",x"4f",x"7f",x"47",x"7f",x"7f",x"7f",x"ed",x"4f",x"df",x"d0",x"4f",x"4f",x"5f",x"6f",x"3f",x"45",x"04",x"20",x"24",x"0f",x"16",x"40",x"10",x"1f",x"2f",x"03",x"2d",x"10",x"11",x"00",x"01",x"28",x"07",x"40",x"10",x"12",x"21",x"1f",x"e2",x"00",x"72",x"34",x"40",x"02",x"00",x"13",x"00",x"02",x"2f",x"f3",x"ad",x"10",x"28",x"30",x"04",x"1f",x"1f",x"2f",x"2f",x"0d",x"10",x"80",x"10",x"44",x"16",x"6f",x"1f",x"2f",x"3f",x"00",x"03",x"2d",x"10",x"10",x"ad",x"10",x"b8",x"13",x"d7",x"cf",x"1f",x"6d",x"10",x"00",x"03",x"ad",x"10",x"ed",x"10",x"03",x"16",x"1f",x"1f",x"2f",x"2f",x"0d",x"10",x"2c",x"20",x"1f",x"f6",x"80",x"10",x"38",x"80",x"10",x"00",x"1f",x"18",x"16",x"18",x"20",x"10",x"28",x"30",x"00",x"1f",x"2f",x"03",x"ed",x"10",x"11",x"00",x"01",x"20",x"04",x"28",x"30",x"0b",x"11",x"40",x"10",x"2f",x"21",x"21",x"60",x"10",x"10",x"30",x"28",x"80",x"04",x"20",x"2c",x"24",x"1a",x"c6",x"7f",x"04",x"28",x"4d",x"10",x"20",x"1f",x"62",x"ff",x"ff",x"1f",x"1f",x"2f",x"7f",x"2f",x"18",x"10",x"28",x"30",x"10",x"28",x"30",x"1f",x"18",x"2f",x"7f",x"35",x"40",x"10",x"2f",x"32",x"80",x"10",x"07",x"2c",x"7f",x"a0",x"10",x"44",x"18",x"28",x"00",x"1f",x"42",x"80",x"04",x"ad",x"10",x"18",x"2d",x"10",x"24",x"1f",x"2f",x"6d",x"10",x"20",x"68",x"18",x"e0",x"10",x"28",x"c0",x"10",x"2c",x"60",x"10",x"10",x"9f",x"08",x"73",x"51",x"1f",x"40",x"02",x"a0",x"1f",x"02",x"4f",x"10",x"ff",x"73",x"f3",x"77",x"00",x"10",x"13",x"00",x"c0",x"23",x"75",x"75",x"ff",x"1a",x"00",x"8a",x"80",x"02",x"6f",x"5f",x"4f",x"df",x"d0",x"00",x"17",x"4f",x"7f",x"7f",x"7f",x"7f",x"7f",x"cd",x"10",x"10",x"4f",x"10",x"cf",x"63",x"4f",x"0f",x"7f",x"7f",x"7f",x"cd",x"10",x"10",x"4f",x"10",x"cf",x"1c",x"4f",x"0f",x"7f",x"7f",x"7f",x"cd",x"10",x"10",x"4f",x"10",x"10",x"10",x"10",x"d0",x"00",x"df",x"04",x"16",x"c2",x"83",x"04",x"0f",x"4f",x"df",x"d0",x"00",x"21",x"10",x"21",x"10",x"81",x"07",x"00",x"20",x"17",x"e0",x"10",x"17",x"87",x"09",x"ff",x"40",x"17",x"80",x"10",x"00",x"28",x"08",x"89",x"98",x"00",x"87",x"04",x"08",x"0c",x"07",x"80",x"10",x"10",x"47",x"33",x"ff",x"03",x"00",x"27",x"17",x"40",x"10",x"10",x"17",x"f8",x"df",x"04",x"01",x"78",x"00",x"10",x"80",x"10",x"00",x"ff",x"f7",x"07",x"08",x"08",x"00",x"00",x"f8",x"87",x"73",x"04",x"00",x"48",x"00",x"ed",x"78",x"87",x"28",x"09",x"00",x"87",x"72",x"43",x"13",x"1d",x"c2",x"10",x"23",x"00",x"02",x"02",x"10",x"00",x"17",x"03",x"4f",x"df",x"8f",x"10",x"df",x"0c",x"08",x"f7",x"ff",x"f1",x"04",x"09",x"02",x"08",x"ff",x"f8",x"40",x"10",x"f9",x"40",x"10",x"40",x"10",x"79",x"13",x"08",x"00",x"f1",x"09",x"08",x"ff",x"f8",x"40",x"10",x"f9",x"40",x"10",x"40",x"10",x"91",x"80",x"10",x"18",x"40",x"10",x"19",x"ff",x"40",x"10",x"40",x"10",x"81",x"40",x"10",x"00",x"58",x"8c",x"06",x"11",x"04",x"00",x"08",x"00",x"07",x"00",x"09",x"00",x"98",x"01",x"00",x"00",x"01",x"31",x"e0",x"10",x"ff",x"21",x"58",x"60",x"10",x"02",x"00",x"45",x"32",x"00",x"01",x"40",x"10",x"02",x"00",x"52",x"60",x"10",x"41",x"e0",x"10",x"31",x"e0",x"10",x"01",x"80",x"10",x"04",x"74",x"58",x"a1",x"05",x"11",x"54",x"00",x"08",x"40",x"10",x"40",x"10",x"47",x"40",x"10",x"40",x"10",x"32",x"00",x"a2",x"00",x"3a",x"07",x"14",x"31",x"ff",x"f1",x"12",x"c0",x"10",x"1c",x"00",x"2f",x"08",x"00",x"81",x"81",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"14",x"80",x"71",x"71",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"02",x"18",x"04",x"f5",x"72",x"04",x"18",x"c7",x"09",x"14",x"07",x"20",x"0a",x"00",x"0a",x"00",x"10",x"14",x"18",x"00",x"7f",x"01",x"00",x"12",x"8f",x"96",x"23",x"32",x"04",x"23",x"32",x"10",x"f3",x"55",x"53",x"01",x"32",x"33",x"33",x"07",x"02",x"72",x"04",x"0f",x"f3",x"01",x"13",x"02",x"18",x"10",x"01",x"8f",x"52",x"02",x"23",x"32",x"08",x"23",x"32",x"32",x"aa",x"27",x"73",x"02",x"66",x"32",x"22",x"32",x"23",x"32",x"1e",x"32",x"02",x"23",x"03",x"18",x"04",x"f5",x"6d",x"10",x"c5",x"42",x"11",x"53",x"52",x"a9",x"00",x"03",x"04",x"00",x"46",x"60",x"a9",x"11",x"f5",x"00",x"41",x"9f",x"2f",x"ad",x"10",x"24",x"01",x"28",x"03",x"ad",x"10",x"02",x"02",x"00",x"01",x"24",x"10",x"2f",x"3f",x"32",x"00",x"02",x"32",x"1c",x"14",x"18",x"03",x"1d",x"82",x"00",x"08",x"60",x"10",x"10",x"05",x"04",x"02",x"43",x"c0",x"10",x"1f",x"01",x"12",x"01",x"73",x"13",x"c0",x"10",x"34",x"08",x"21",x"02",x"64",x"40",x"10",x"00",x"40",x"10",x"10",x"80",x"10",x"01",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"18",x"00",x"74",x"48",x"31",x"01",x"54",x"a3",x"8c",x"01",x"51",x"51",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"02",x"18",x"16",x"41",x"63",x"00",x"9f",x"14",x"69",x"f9",x"80",x"10",x"1c",x"ff",x"08",x"21",x"00",x"09",x"00",x"16",x"96",x"21",x"41",x"10",x"ad",x"10",x"01",x"00",x"06",x"10",x"52",x"0f",x"14",x"05",x"41",x"ff",x"f2",x"03",x"18",x"41",x"31",x"31",x"1c",x"93",x"32",x"53",x"40",x"10",x"18",x"01",x"c0",x"10",x"03",x"28",x"8c",x"04",x"08",x"0c",x"cf",x"10",x"37",x"20",x"10",x"e0",x"12",x"02",x"10",x"a0",x"10",x"31",x"37",x"72",x"32",x"03",x"31",x"d0",x"00",x"17",x"4f",x"40",x"10",x"ff",x"f9",x"91",x"00",x"08",x"00",x"0b",x"00",x"ba",x"0a",x"00",x"39",x"1b",x"40",x"10",x"1e",x"ff",x"40",x"10",x"40",x"10",x"ba",x"60",x"10",x"07",x"08",x"07",x"20",x"10",x"07",x"60",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"80",x"10",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"40",x"10",x"78",x"08",x"00",x"17",x"42",x"01",x"00",x"07",x"71",x"d0",x"00",x"17",x"4f",x"40",x"10",x"ff",x"f9",x"91",x"00",x"08",x"00",x"0b",x"00",x"ba",x"f7",x"80",x"10",x"1a",x"04",x"00",x"0b",x"00",x"09",x"00",x"0e",x"00",x"eb",x"0a",x"00",x"89",x"24",x"78",x"08",x"00",x"13",x"07",x"00",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"20",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"98",x"07",x"40",x"10",x"31",x"21",x"40",x"10",x"4f",x"4f",x"10",x"ff",x"f7",x"12",x"17",x"40",x"10",x"00",x"07",x"40",x"10",x"40",x"10",x"12",x"e0",x"10",x"ff",x"12",x"13",x"40",x"10",x"00",x"03",x"00",x"02",x"00",x"21",x"4f",x"10",x"cf",x"1a",x"02",x"00",x"0a",x"ff",x"1b",x"08",x"ff",x"40",x"10",x"40",x"10",x"7a",x"80",x"10",x"1a",x"04",x"00",x"0b",x"00",x"09",x"00",x"0e",x"00",x"eb",x"0a",x"00",x"89",x"24",x"78",x"08",x"00",x"13",x"07",x"00",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"20",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"98",x"f7",x"40",x"10",x"31",x"21",x"40",x"10",x"4f",x"4f",x"10",x"cf",x"1a",x"02",x"00",x"0a",x"ff",x"1b",x"08",x"ff",x"40",x"10",x"40",x"10",x"7a",x"80",x"10",x"1a",x"04",x"00",x"0b",x"00",x"09",x"00",x"0e",x"00",x"eb",x"0a",x"00",x"89",x"24",x"78",x"08",x"00",x"13",x"07",x"00",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"20",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"98",x"f7",x"40",x"10",x"31",x"21",x"40",x"10",x"4f",x"4f",x"10",x"cf",x"1a",x"02",x"00",x"0a",x"ff",x"1b",x"08",x"ff",x"40",x"10",x"40",x"10",x"7a",x"80",x"10",x"1a",x"04",x"00",x"0b",x"00",x"09",x"00",x"0e",x"00",x"eb",x"0a",x"00",x"89",x"24",x"78",x"08",x"00",x"13",x"07",x"00",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"20",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"98",x"f7",x"40",x"10",x"31",x"21",x"40",x"10",x"4f",x"4f",x"10",x"cf",x"1a",x"02",x"00",x"0a",x"ff",x"1b",x"08",x"ff",x"40",x"10",x"40",x"10",x"7a",x"0a",x"00",x"39",x"1b",x"40",x"10",x"1e",x"ff",x"40",x"10",x"40",x"10",x"ba",x"60",x"10",x"07",x"08",x"07",x"20",x"10",x"07",x"60",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"80",x"10",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"40",x"10",x"87",x"f7",x"00",x"17",x"42",x"01",x"00",x"07",x"71",x"d0",x"00",x"2e",x"02",x"00",x"df",x"0c",x"08",x"04",x"37",x"2f",x"f2",x"27",x"28",x"14",x"ff",x"f2",x"08",x"7f",x"2f",x"72",x"d2",x"80",x"10",x"28",x"e2",x"80",x"10",x"00",x"ff",x"f7",x"10",x"19",x"71",x"40",x"10",x"1a",x"ff",x"40",x"10",x"40",x"10",x"98",x"20",x"10",x"00",x"21",x"a0",x"10",x"05",x"17",x"40",x"10",x"18",x"ff",x"40",x"10",x"9f",x"40",x"10",x"71",x"00",x"10",x"00",x"4e",x"09",x"03",x"01",x"10",x"20",x"00",x"4f",x"42",x"03",x"1f",x"11",x"12",x"f3",x"31",x"06",x"45",x"30",x"6d",x"10",x"03",x"12",x"01",x"0d",x"c2",x"11",x"03",x"12",x"01",x"ad",x"10",x"03",x"12",x"01",x"0d",x"c2",x"11",x"03",x"12",x"01",x"ed",x"10",x"03",x"12",x"01",x"0d",x"c2",x"11",x"03",x"16",x"1f",x"62",x"0b",x"ad",x"10",x"30",x"01",x"03",x"0c",x"5c",x"02",x"64",x"02",x"03",x"01",x"0c",x"1f",x"01",x"03",x"ad",x"10",x"30",x"f7",x"31",x"32",x"05",x"30",x"38",x"14",x"10",x"02",x"1e",x"00",x"03",x"04",x"03",x"0c",x"1f",x"01",x"03",x"14",x"0c",x"2f",x"64",x"03",x"05",x"21",x"2f",x"01",x"0c",x"15",x"03",x"1f",x"c1",x"30",x"06",x"6d",x"10",x"14",x"03",x"02",x"32",x"02",x"03",x"34",x"05",x"28",x"2c",x"00",x"12",x"2f",x"12",x"20",x"10",x"14",x"51",x"1c",x"18",x"0b",x"2f",x"03",x"c3",x"15",x"80",x"00",x"01",x"03",x"03",x"00",x"51",x"01",x"01",x"60",x"10",x"1f",x"01",x"01",x"51",x"14",x"1c",x"18",x"0b",x"2f",x"03",x"22",x"12",x"24",x"00",x"f1",x"80",x"10",x"01",x"bf",x"01",x"00",x"60",x"af",x"33",x"22",x"02",x"13",x"00",x"03",x"40",x"10",x"40",x"10",x"ff",x"f7",x"14",x"71",x"14",x"21",x"23",x"19",x"00",x"51",x"01",x"00",x"0e",x"00",x"0e",x"00",x"7f",x"2e",x"01",x"00",x"80",x"10",x"01",x"e0",x"10",x"ff",x"f2",x"01",x"07",x"00",x"71",x"71",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"16",x"80",x"10",x"ff",x"0e",x"c0",x"54",x"01",x"00",x"0e",x"10",x"ff",x"0e",x"04",x"08",x"0c",x"91",x"cf",x"10",x"01",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"11",x"21",x"63",x"71",x"ad",x"10",x"c1",x"61",x"8f",x"ff",x"f5",x"00",x"60",x"ef",x"08",x"00",x"81",x"7f",x"81",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"15",x"e0",x"7f",x"ef",x"6f",x"e0",x"10",x"01",x"14",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"11",x"21",x"53",x"81",x"ed",x"10",x"56",x"c4",x"1f",x"20",x"10",x"df",x"08",x"04",x"24",x"1f",x"02",x"01",x"1f",x"03",x"02",x"08",x"45",x"5f",x"4f",x"df",x"1f",x"21",x"cf",x"10",x"df",x"04",x"f4",x"40",x"10",x"ff",x"f1",x"00",x"31",x"14",x"f7",x"73",x"ff",x"37",x"00",x"43",x"03",x"01",x"60",x"03",x"60",x"10",x"cc",x"f2",x"c2",x"07",x"c3",x"04",x"31",x"d0",x"00",x"14",x"07",x"03",x"ff",x"08",x"00",x"01",x"00",x"22",x"11",x"e3",x"21",x"00",x"73",x"21",x"03",x"d0",x"00",x"12",x"03",x"4f",x"02",x"00",x"21",x"21",x"02",x"13",x"31",x"08",x"13",x"31",x"31",x"aa",x"17",x"73",x"01",x"66",x"31",x"11",x"31",x"13",x"31",x"1e",x"31",x"02",x"13",x"f3",x"18",x"04",x"41",x"01",x"f1",x"00",x"02",x"21",x"14",x"00",x"01",x"04",x"3c",x"d0",x"00",x"37",x"00",x"10",x"e0",x"02",x"e0",x"03",x"00",x"07",x"02",x"07",x"07",x"01",x"03",x"2c",x"10",x"df",x"08",x"04",x"14",x"fd",x"15",x"5f",x"14",x"4f",x"df",x"d0",x"00",x"df",x"0c",x"08",x"04",x"31",x"00",x"07",x"72",x"14",x"10",x"07",x"7f",x"17",x"27",x"00",x"23",x"12",x"24",x"18",x"14",x"ff",x"07",x"00",x"2f",x"f2",x"07",x"00",x"00",x"10",x"ff",x"18",x"06",x"02",x"00",x"09",x"00",x"02",x"00",x"0a",x"00",x"a9",x"08",x"00",x"00",x"02",x"03",x"03",x"73",x"11",x"0b",x"00",x"07",x"00",x"04",x"00",x"08",x"00",x"87",x"01",x"01",x"00",x"01",x"13",x"03",x"01",x"1c",x"0b",x"03",x"6f",x"b6",x"ed",x"10",x"30",x"28",x"15",x"1f",x"11",x"12",x"1f",x"00",x"02",x"04",x"52",x"18",x"04",x"1f",x"00",x"01",x"2f",x"16",x"01",x"c1",x"06",x"52",x"1f",x"01",x"2c",x"04",x"1f",x"c6",x"03",x"30",x"52",x"30",x"4f",x"2d",x"10",x"14",x"2c",x"c2",x"72",x"30",x"03",x"08",x"f8",x"09",x"00",x"19",x"1f",x"07",x"1f",x"3f",x"31",x"1c",x"11",x"00",x"10",x"c0",x"00",x"01",x"03",x"03",x"00",x"3f",x"4b",x"01",x"00",x"80",x"88",x"63",x"37",x"99",x"66",x"10",x"f1",x"60",x"10",x"10",x"60",x"10",x"10",x"14",x"00",x"11",x"92",x"40",x"10",x"10",x"b1",x"00",x"10",x"01",x"20",x"10",x"ff",x"06",x"c0",x"10",x"ff",x"06",x"01",x"17",x"1c",x"18",x"05",x"05",x"14",x"00",x"06",x"01",x"7f",x"26",x"01",x"00",x"c0",x"10",x"01",x"80",x"10",x"01",x"05",x"00",x"20",x"10",x"40",x"10",x"01",x"1c",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"18",x"01",x"a1",x"26",x"ad",x"10",x"1f",x"41",x"24",x"03",x"3f",x"6d",x"10",x"01",x"00",x"01",x"14",x"1c",x"18",x"28",x"62",x"ec",x"2f",x"53",x"1f",x"1f",x"2f",x"c1",x"62",x"14",x"2d",x"10",x"20",x"02",x"17",x"00",x"40",x"10",x"9f",x"09",x"00",x"03",x"00",x"73",x"10",x"07",x"73",x"21",x"00",x"01",x"91",x"80",x"10",x"02",x"16",x"a0",x"06",x"10",x"6c",x"04",x"08",x"0c",x"31",x"d0",x"61",x"bf",x"61",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"02",x"18",x"05",x"f5",x"62",x"eb",x"bf",x"17",x"c6",x"05",x"00",x"60",x"10",x"10",x"18",x"80",x"10",x"01",x"14",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"18",x"10",x"14",x"1c",x"fb",x"b1",x"7f",x"b1",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"02",x"18",x"04",x"f5",x"b2",x"ea",x"1f",x"51",x"cb",x"01",x"1c",x"fa",x"00",x"29",x"48",x"14",x"4f",x"07",x"ff",x"f1",x"0a",x"0b",x"ab",x"a9",x"ea",x"a9",x"0a",x"02",x"03",x"08",x"a7",x"10",x"83",x"10",x"10",x"3c",x"4f",x"10",x"00",x"07",x"4f",x"73",x"e2",x"4f",x"df",x"d0",x"00",x"02",x"01",x"01",x"01",x"17",x"17",x"02",x"78",x"87",x"08",x"28",x"82",x"78",x"78",x"02",x"79",x"79",x"87",x"55",x"58",x"01",x"ba",x"9b",x"b9",x"10",x"33",x"39",x"9a",x"aa",x"9a",x"01",x"ea",x"08",x"04",x"98",x"88",x"98",x"89",x"98",x"1e",x"98",x"01",x"19",x"07",x"08",x"18",x"18",x"08",x"40",x"10",x"00",x"d0",x"f3",x"83",x"18",x"31",x"c0",x"10",x"0a",x"21",x"19",x"1f",x"01",x"01",x"08",x"73",x"0b",x"1f",x"0e",x"07",x"0a",x"ff",x"31",x"17",x"31",x"10",x"df",x"08",x"04",x"14",x"fe",x"15",x"5f",x"14",x"4f",x"df",x"d0",x"00",x"40",x"14",x"52",x"08",x"47",x"bf",x"3a",x"00",x"df",x"e4",x"e9",x"ee",x"bb",x"c4",x"cd",x"d6",x"97",x"a0",x"a9",x"b2",x"73",x"7c",x"85",x"8e",x"74",x"48",x"00",x"63",x"6b",x"72",x"6d",x"65",x"6e",x"72",x"74",x"20",x"20",x"65",x"6b",x"36",x"61",x"61",x"6e",x"6e",x"72",x"74",x"20",x"20",x"65",x"6b",x"50",x"69",x"67",x"72",x"6f",x"75",x"61",x"65",x"73",x"72",x"72",x"72",x"00",x"70",x"6f",x"6e",x"72",x"70",x"6d",x"72",x"6f",x"6f",x"61",x"0a",x"20",x"69",x"69",x"72",x"70",x"6d",x"72",x"6f",x"6f",x"61",x"0a",x"75",x"52",x"20",x"74",x"63",x"25",x"20",x"68",x"64",x"20",x"30",x"00",x"5d",x"4f",x"6d",x"69",x"72",x"78",x"78",x"73",x"6c",x"65",x"25",x"0a",x"75",x"52",x"20",x"74",x"72",x"78",x"78",x"73",x"6c",x"65",x"25",x"0a",x"72",x"72",x"69",x"20",x"20",x"0a",x"74",x"74",x"73",x"20",x"20",x"0a",x"74",x"74",x"20",x"63",x"20",x"00",x"72",x"6f",x"53",x"20",x"25",x"45",x"52",x"75",x"65",x"75",x"66",x"61",x"65",x"20",x"73",x"20",x"20",x"61",x"20",x"75",x"0a",x"65",x"69",x"20",x"20",x"20",x"0a",x"6d",x"65",x"65",x"6f",x"20",x"00",x"34",x"31",x"6d",x"69",x"20",x"6e",x"2e",x"74",x"2f",x"45",x"5f",x"66",x"6c",x"6f",x"6c",x"66",x"73",x"3a",x"0a",x"6d",x"20",x"61",x"6e",x"20",x"00",x"43",x"65",x"72",x"20",x"20",x"3a",x"25",x"0a",x"64",x"63",x"74",x"20",x"3a",x"25",x"0a",x"64",x"63",x"72",x"20",x"3a",x"25",x"0a",x"64",x"63",x"74",x"20",x"3a",x"25",x"0a",x"64",x"63",x"61",x"20",x"3a",x"25",x"0a",x"72",x"74",x"65",x"69",x"76",x"64",x"64",x"65",x"65",x"65",x"74",x"72",x"6e",x"64",x"70",x"69",x"72",x"73",x"43",x"4d",x"20",x"20",x"66",x"25",x"73",x"20",x"45",x"72",x"65",x"74",x"00",x"6e",x"76",x"64",x"20",x"72",x"6f",x"6f",x"68",x"20",x"64",x"6c",x"2c",x"65",x"20",x"70",x"20",x"68",x"73",x"73",x"20",x"6e",x"20",x"74",x"6d",x"54",x"65",x"00",x"54",x"71",x"33",x"34",x"34",x"2d",x"35",x"30",x"00",x"32",x"32",x"37",x"33",x"30",x"2d",x"33",x"34",x"00",x"33",x"30",x"31",x"30",x"30",x"34",x"35",x"00",x"34",x"37",x"31",x"3c",x"4c",x"31",x"35",x"39",x"64",x"68",x"6c",x"70",x"74",x"78",x"30",x"34",x"38",x"43",x"47",x"4b",x"4f",x"53",x"57",x"00",x"00",x"50",x"57",x"5c",x"00",x"66",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
 shared variable RAM1: RAM_TABLE := RAM_TABLE'(
x"60",x"18",x"70",x"fe",x"70",x"40",x"70",x"10",x"60",x"98",x"18",x"40",x"38",x"40",x"40",x"70",x"70",x"18",x"07",x"50",x"46",x"00",x"00",x"00",x"f4",x"70",x"38",x"40",x"cf",x"20",x"24",x"30",x"4f",x"4f",x"00",x"10",x"40",x"40",x"40",x"40",x"19",x"f8",x"04",x"c0",x"38",x"04",x"40",x"89",x"70",x"88",x"05",x"04",x"c0",x"38",x"38",x"40",x"98",x"98",x"99",x"19",x"40",x"40",x"c0",x"38",x"3a",x"0c",x"40",x"40",x"0c",x"40",x"40",x"c4",x"38",x"40",x"38",x"c0",x"38",x"38",x"40",x"40",x"40",x"40",x"0c",x"40",x"40",x"c1",x"38",x"40",x"38",x"40",x"40",x"19",x"60",x"04",x"40",x"11",x"60",x"f8",x"98",x"04",x"04",x"05",x"40",x"98",x"98",x"98",x"18",x"30",x"00",x"10",x"40",x"90",x"0c",x"40",x"cb",x"38",x"0c",x"cb",x"38",x"20",x"40",x"40",x"40",x"51",x"38",x"c2",x"38",x"3a",x"60",x"84",x"89",x"ff",x"04",x"11",x"3a",x"89",x"04",x"11",x"40",x"40",x"3a",x"20",x"38",x"11",x"40",x"40",x"38",x"10",x"40",x"40",x"40",x"40",x"40",x"40",x"70",x"90",x"c0",x"38",x"40",x"80",x"00",x"80",x"7f",x"ff",x"70",x"90",x"70",x"40",x"90",x"0c",x"6f",x"43",x"42",x"98",x"84",x"99",x"07",x"41",x"43",x"18",x"60",x"42",x"4d",x"84",x"0c",x"40",x"40",x"c0",x"38",x"38",x"70",x"ce",x"38",x"38",x"40",x"0c",x"60",x"42",x"0c",x"10",x"60",x"41",x"0c",x"c1",x"38",x"50",x"40",x"98",x"04",x"90",x"43",x"98",x"19",x"84",x"60",x"42",x"98",x"89",x"04",x"00",x"40",x"50",x"c0",x"38",x"10",x"10",x"80",x"70",x"04",x"40",x"00",x"07",x"45",x"98",x"ff",x"04",x"40",x"40",x"38",x"70",x"0c",x"40",x"40",x"82",x"c1",x"38",x"40",x"fb",x"ce",x"38",x"98",x"00",x"18",x"40",x"40",x"40",x"40",x"40",x"18",x"3a",x"6f",x"43",x"43",x"60",x"42",x"80",x"7f",x"0c",x"40",x"40",x"c4",x"38",x"60",x"41",x"42",x"98",x"60",x"42",x"0c",x"40",x"40",x"c1",x"38",x"60",x"41",x"18",x"c2",x"38",x"60",x"84",x"98",x"19",x"c8",x"38",x"0c",x"cd",x"38",x"40",x"98",x"98",x"90",x"90",x"70",x"10",x"0c",x"40",x"40",x"0c",x"60",x"42",x"80",x"7f",x"20",x"40",x"3a",x"40",x"18",x"60",x"41",x"80",x"7f",x"40",x"40",x"98",x"18",x"30",x"0c",x"40",x"70",x"c0",x"38",x"38",x"c5",x"38",x"60",x"04",x"40",x"40",x"c0",x"38",x"38",x"60",x"41",x"42",x"60",x"42",x"19",x"98",x"9a",x"07",x"41",x"41",x"18",x"ce",x"38",x"38",x"30",x"0c",x"38",x"60",x"41",x"41",x"0c",x"10",x"60",x"41",x"0c",x"38",x"0c",x"38",x"0c",x"10",x"40",x"40",x"40",x"40",x"40",x"40",x"c0",x"38",x"40",x"70",x"70",x"0c",x"50",x"40",x"98",x"90",x"70",x"40",x"0c",x"46",x"cf",x"38",x"0c",x"40",x"c2",x"38",x"c4",x"38",x"c4",x"38",x"c1",x"38",x"5f",x"0c",x"41",x"60",x"42",x"60",x"41",x"18",x"0c",x"98",x"60",x"41",x"47",x"10",x"38",x"40",x"cb",x"38",x"0c",x"90",x"98",x"60",x"c8",x"38",x"38",x"40",x"0c",x"98",x"98",x"98",x"98",x"30",x"60",x"43",x"98",x"18",x"0c",x"5f",x"38",x"98",x"0c",x"0c",x"c7",x"38",x"40",x"40",x"98",x"98",x"0c",x"18",x"60",x"41",x"41",x"98",x"07",x"45",x"90",x"40",x"90",x"70",x"40",x"98",x"ce",x"38",x"40",x"10",x"40",x"40",x"40",x"40",x"c7",x"38",x"40",x"40",x"40",x"52",x"38",x"40",x"18",x"40",x"40",x"40",x"40",x"18",x"0c",x"30",x"98",x"98",x"90",x"90",x"18",x"10",x"38",x"5e",x"90",x"0c",x"90",x"90",x"90",x"ca",x"38",x"40",x"10",x"40",x"88",x"80",x"80",x"90",x"91",x"80",x"78",x"88",x"80",x"c4",x"38",x"40",x"40",x"c4",x"38",x"80",x"70",x"40",x"ff",x"90",x"91",x"80",x"7f",x"0c",x"40",x"20",x"41",x"60",x"40",x"42",x"98",x"80",x"7f",x"04",x"40",x"c4",x"38",x"40",x"c3",x"38",x"70",x"84",x"86",x"88",x"04",x"20",x"40",x"20",x"0c",x"ff",x"10",x"40",x"11",x"40",x"98",x"50",x"ca",x"38",x"18",x"c5",x"38",x"40",x"40",x"60",x"84",x"70",x"40",x"70",x"40",x"40",x"40",x"c0",x"38",x"40",x"04",x"05",x"40",x"40",x"18",x"0c",x"41",x"0c",x"40",x"c8",x"38",x"40",x"40",x"40",x"51",x"38",x"90",x"98",x"70",x"80",x"07",x"48",x"18",x"40",x"07",x"48",x"10",x"18",x"10",x"90",x"18",x"10",x"40",x"11",x"40",x"40",x"40",x"50",x"38",x"10",x"40",x"90",x"90",x"70",x"40",x"40",x"40",x"40",x"40",x"c4",x"38",x"70",x"40",x"99",x"ca",x"38",x"40",x"7f",x"40",x"99",x"c8",x"38",x"40",x"c0",x"38",x"40",x"07",x"49",x"98",x"98",x"98",x"18",x"51",x"38",x"d9",x"10",x"40",x"40",x"40",x"40",x"40",x"8c",x"80",x"90",x"54",x"60",x"40",x"40",x"70",x"40",x"91",x"70",x"40",x"91",x"70",x"40",x"91",x"70",x"40",x"90",x"70",x"40",x"70",x"c0",x"38",x"90",x"99",x"60",x"42",x"43",x"99",x"70",x"c6",x"38",x"40",x"60",x"41",x"f1",x"76",x"40",x"40",x"40",x"40",x"38",x"c2",x"38",x"40",x"60",x"41",x"99",x"60",x"41",x"70",x"91",x"91",x"91",x"99",x"8c",x"70",x"60",x"40",x"40",x"40",x"40",x"70",x"20",x"04",x"80",x"90",x"89",x"91",x"90",x"80",x"90",x"89",x"80",x"90",x"00",x"80",x"7f",x"fd",x"ce",x"38",x"60",x"40",x"90",x"60",x"42",x"70",x"40",x"60",x"40",x"c1",x"38",x"82",x"50",x"00",x"40",x"60",x"40",x"60",x"40",x"c1",x"38",x"60",x"04",x"20",x"90",x"60",x"42",x"98",x"3a",x"40",x"90",x"98",x"70",x"60",x"42",x"99",x"99",x"88",x"3a",x"20",x"60",x"40",x"40",x"40",x"40",x"40",x"98",x"70",x"60",x"42",x"99",x"98",x"3a",x"40",x"40",x"98",x"60",x"41",x"70",x"40",x"40",x"98",x"70",x"20",x"40",x"40",x"8c",x"cf",x"38",x"40",x"cf",x"38",x"40",x"0c",x"60",x"70",x"60",x"40",x"ce",x"38",x"60",x"41",x"70",x"60",x"40",x"f0",x"70",x"cc",x"38",x"70",x"43",x"70",x"70",x"60",x"41",x"c7",x"38",x"60",x"40",x"c4",x"38",x"60",x"42",x"0c",x"c4",x"38",x"40",x"8b",x"90",x"c5",x"38",x"40",x"60",x"40",x"40",x"c4",x"38",x"40",x"0c",x"40",x"3a",x"40",x"0c",x"40",x"c8",x"38",x"99",x"3a",x"40",x"0c",x"40",x"c6",x"38",x"80",x"7f",x"e0",x"c2",x"38",x"40",x"42",x"43",x"f1",x"cb",x"38",x"46",x"e0",x"c3",x"38",x"60",x"c0",x"38",x"38",x"40",x"40",x"70",x"38",x"40",x"41",x"fb",x"c6",x"38",x"42",x"f8",x"c5",x"38",x"41",x"80",x"60",x"41",x"f6",x"c4",x"38",x"f6",x"70",x"60",x"42",x"80",x"90",x"80",x"90",x"88",x"80",x"90",x"ff",x"70",x"00",x"60",x"40",x"40",x"80",x"90",x"f0",x"00",x"80",x"90",x"80",x"90",x"80",x"90",x"74",x"60",x"40",x"20",x"20",x"91",x"70",x"40",x"60",x"41",x"70",x"38",x"40",x"60",x"40",x"70",x"c1",x"38",x"40",x"c8",x"38",x"40",x"91",x"98",x"70",x"60",x"42",x"99",x"80",x"98",x"19",x"c1",x"38",x"40",x"c4",x"38",x"40",x"91",x"98",x"70",x"60",x"42",x"99",x"80",x"98",x"19",x"c1",x"38",x"40",x"c0",x"38",x"40",x"91",x"80",x"98",x"80",x"98",x"00",x"80",x"7f",x"20",x"40",x"07",x"49",x"80",x"98",x"80",x"98",x"80",x"98",x"80",x"90",x"80",x"90",x"80",x"90",x"80",x"90",x"c5",x"38",x"60",x"40",x"40",x"40",x"40",x"fe",x"0c",x"40",x"0c",x"40",x"0c",x"40",x"c5",x"38",x"c8",x"38",x"70",x"0c",x"60",x"40",x"40",x"70",x"c0",x"38",x"80",x"98",x"0c",x"70",x"40",x"60",x"c0",x"38",x"05",x"60",x"40",x"04",x"c3",x"38",x"40",x"40",x"8b",x"c2",x"38",x"0c",x"c1",x"38",x"0c",x"0c",x"40",x"0c",x"40",x"cc",x"38",x"ce",x"38",x"a4",x"70",x"0c",x"60",x"40",x"40",x"70",x"c0",x"38",x"80",x"98",x"0c",x"60",x"70",x"40",x"6f",x"c0",x"38",x"80",x"98",x"80",x"98",x"80",x"98",x"05",x"20",x"04",x"c0",x"38",x"40",x"40",x"50",x"40",x"40",x"8b",x"f7",x"c2",x"38",x"40",x"40",x"40",x"fd",x"f7",x"c0",x"38",x"40",x"40",x"40",x"f0",x"0c",x"40",x"98",x"70",x"60",x"41",x"80",x"90",x"45",x"80",x"90",x"18",x"c4",x"38",x"60",x"40",x"f6",x"70",x"8b",x"00",x"40",x"40",x"40",x"50",x"60",x"84",x"18",x"cd",x"38",x"40",x"40",x"04",x"c4",x"38",x"60",x"42",x"80",x"98",x"70",x"40",x"74",x"20",x"99",x"f4",x"c3",x"38",x"80",x"7f",x"20",x"07",x"49",x"98",x"70",x"f6",x"60",x"80",x"98",x"c4",x"38",x"c7",x"38",x"f6",x"70",x"0c",x"20",x"99",x"f5",x"ce",x"38",x"80",x"7f",x"84",x"18",x"cd",x"38",x"c3",x"38",x"f6",x"70",x"0c",x"20",x"99",x"f7",x"ca",x"38",x"80",x"7f",x"84",x"18",x"cd",x"38",x"60",x"40",x"60",x"04",x"c0",x"38",x"38",x"60",x"45",x"ff",x"c8",x"38",x"40",x"40",x"80",x"98",x"60",x"41",x"f6",x"98",x"18",x"20",x"40",x"0c",x"60",x"40",x"c4",x"38",x"0c",x"0c",x"40",x"0c",x"40",x"fa",x"90",x"fd",x"cf",x"38",x"40",x"40",x"40",x"f6",x"40",x"f1",x"cd",x"38",x"60",x"40",x"40",x"98",x"98",x"98",x"18",x"d6",x"30",x"00",x"10",x"40",x"40",x"98",x"98",x"98",x"18",x"40",x"41",x"0c",x"40",x"98",x"98",x"18",x"30",x"5d",x"40",x"90",x"90",x"0c",x"90",x"60",x"42",x"f0",x"05",x"40",x"8b",x"70",x"20",x"07",x"40",x"19",x"11",x"49",x"50",x"cd",x"38",x"8b",x"70",x"20",x"07",x"40",x"40",x"00",x"3a",x"20",x"cd",x"38",x"07",x"49",x"90",x"70",x"70",x"8b",x"70",x"20",x"40",x"18",x"40",x"07",x"46",x"50",x"41",x"70",x"c0",x"38",x"00",x"0c",x"cc",x"38",x"0c",x"cb",x"38",x"70",x"c0",x"38",x"40",x"70",x"88",x"8b",x"70",x"00",x"80",x"88",x"50",x"88",x"00",x"19",x"3a",x"8b",x"00",x"49",x"50",x"07",x"49",x"70",x"70",x"8b",x"70",x"20",x"40",x"18",x"40",x"07",x"46",x"50",x"41",x"0c",x"07",x"43",x"70",x"0c",x"0c",x"cc",x"38",x"0c",x"cb",x"38",x"0c",x"40",x"0c",x"ce",x"38",x"40",x"0c",x"40",x"20",x"80",x"0c",x"70",x"40",x"10",x"20",x"20",x"07",x"88",x"88",x"00",x"19",x"3a",x"8b",x"00",x"49",x"50",x"10",x"cb",x"38",x"07",x"49",x"98",x"70",x"70",x"8b",x"70",x"20",x"40",x"18",x"07",x"46",x"50",x"41",x"0c",x"07",x"43",x"70",x"0c",x"0c",x"cc",x"38",x"0c",x"cb",x"38",x"40",x"0c",x"40",x"0c",x"c5",x"38",x"90",x"70",x"70",x"40",x"40",x"20",x"90",x"80",x"70",x"40",x"20",x"10",x"20",x"40",x"19",x"8b",x"50",x"00",x"40",x"19",x"8b",x"89",x"89",x"04",x"8b",x"00",x"49",x"10",x"98",x"07",x"49",x"98",x"50",x"c8",x"38",x"70",x"70",x"20",x"80",x"88",x"00",x"98",x"00",x"c0",x"38",x"70",x"38",x"07",x"43",x"70",x"50",x"07",x"49",x"50",x"07",x"49",x"98",x"42",x"70",x"90",x"c7",x"38",x"70",x"40",x"0c",x"70",x"40",x"0c",x"c5",x"38",x"c4",x"38",x"40",x"40",x"8b",x"70",x"20",x"07",x"40",x"19",x"20",x"ce",x"38",x"07",x"49",x"40",x"70",x"40",x"98",x"98",x"98",x"18",x"52",x"38",x"c2",x"38",x"8b",x"70",x"20",x"07",x"40",x"19",x"11",x"49",x"50",x"cd",x"38",x"38",x"5f",x"60",x"42",x"70",x"20",x"80",x"50",x"88",x"88",x"00",x"19",x"8b",x"10",x"49",x"50",x"cc",x"38",x"50",x"38",x"70",x"40",x"60",x"42",x"70",x"70",x"8b",x"70",x"20",x"40",x"18",x"07",x"46",x"50",x"41",x"70",x"c0",x"38",x"00",x"0c",x"cc",x"38",x"0c",x"cb",x"38",x"98",x"3a",x"30",x"5f",x"40",x"60",x"42",x"70",x"40",x"20",x"70",x"10",x"20",x"40",x"07",x"40",x"00",x"19",x"3a",x"20",x"cd",x"38",x"10",x"cb",x"38",x"98",x"50",x"38",x"90",x"90",x"10",x"c5",x"38",x"8b",x"70",x"20",x"70",x"40",x"10",x"20",x"20",x"07",x"88",x"88",x"00",x"19",x"3a",x"8b",x"00",x"49",x"50",x"07",x"49",x"50",x"ca",x"38",x"98",x"98",x"50",x"38",x"90",x"90",x"10",x"40",x"c8",x"38",x"77",x"8b",x"70",x"40",x"40",x"20",x"70",x"40",x"20",x"8b",x"80",x"50",x"00",x"40",x"40",x"00",x"19",x"3a",x"20",x"40",x"40",x"04",x"20",x"cc",x"38",x"10",x"ca",x"38",x"40",x"07",x"49",x"18",x"40",x"40",x"30",x"00",x"0c",x"90",x"90",x"10",x"40",x"c0",x"38",x"7f",x"c1",x"38",x"0c",x"40",x"20",x"40",x"ce",x"38",x"7f",x"04",x"20",x"42",x"70",x"8b",x"70",x"8b",x"ff",x"70",x"40",x"40",x"04",x"20",x"20",x"07",x"20",x"40",x"40",x"80",x"80",x"11",x"ff",x"50",x"11",x"49",x"50",x"07",x"49",x"98",x"88",x"88",x"00",x"40",x"90",x"90",x"10",x"98",x"98",x"51",x"38",x"10",x"40",x"40",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"0c",x"90",x"1a",x"c0",x"38",x"38",x"40",x"40",x"40",x"88",x"8c",x"00",x"50",x"98",x"1a",x"c0",x"38",x"38",x"40",x"90",x"60",x"20",x"40",x"45",x"0c",x"62",x"42",x"06",x"00",x"ce",x"38",x"40",x"40",x"1a",x"c0",x"38",x"38",x"40",x"40",x"40",x"88",x"8c",x"00",x"50",x"98",x"1a",x"c0",x"38",x"38",x"40",x"40",x"c2",x"38",x"40",x"62",x"42",x"06",x"00",x"ce",x"38",x"40",x"40",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"0c",x"40",x"40",x"98",x"98",x"98",x"18",x"30",x"00",x"70",x"60",x"41",x"cd",x"38",x"ff",x"72",x"20",x"c0",x"38",x"40",x"60",x"47",x"60",x"42",x"60",x"42",x"cb",x"38",x"40",x"60",x"47",x"98",x"50",x"40",x"c5",x"38",x"c2",x"38",x"c0",x"38",x"40",x"62",x"41",x"98",x"50",x"40",x"c2",x"38",x"c0",x"38",x"40",x"98",x"50",x"40",x"40",x"20",x"60",x"49",x"cb",x"38",x"40",x"20",x"60",x"49",x"70",x"cd",x"38",x"cd",x"38",x"cc",x"38",x"cc",x"38",x"cc",x"38",x"c0",x"38",x"ce",x"38",x"40",x"90",x"70",x"40",x"60",x"41",x"85",x"04",x"c6",x"38",x"40",x"90",x"70",x"38",x"c7",x"38",x"40",x"20",x"60",x"49",x"c9",x"38",x"40",x"50",x"40",x"c4",x"38",x"44",x"80",x"84",x"70",x"c2",x"38",x"38",x"40",x"20",x"60",x"49",x"46",x"98",x"50",x"40",x"18",x"10",x"40",x"40",x"c1",x"38",x"60",x"41",x"40",x"0c",x"38",x"40",x"0c",x"38",x"40",x"90",x"42",x"98",x"50",x"40",x"38",x"40",x"90",x"40",x"98",x"50",x"40",x"40",x"4b",x"5e",x"90",x"90",x"90",x"90",x"80",x"70",x"70",x"40",x"80",x"70",x"70",x"20",x"20",x"40",x"c0",x"38",x"40",x"70",x"c2",x"38",x"20",x"20",x"07",x"1a",x"ce",x"38",x"80",x"12",x"70",x"84",x"60",x"47",x"60",x"49",x"80",x"60",x"48",x"45",x"80",x"60",x"49",x"60",x"41",x"89",x"70",x"f4",x"c6",x"38",x"40",x"04",x"40",x"40",x"89",x"70",x"f1",x"80",x"70",x"c4",x"38",x"40",x"04",x"40",x"40",x"98",x"07",x"48",x"80",x"82",x"0c",x"c0",x"38",x"40",x"40",x"40",x"51",x"38",x"70",x"c1",x"38",x"c0",x"38",x"38",x"40",x"38",x"c2",x"38",x"c0",x"38",x"38",x"40",x"38",x"c2",x"38",x"40",x"38",x"40",x"38",x"c0",x"38",x"40",x"30",x"f0",x"86",x"70",x"20",x"c0",x"38",x"89",x"88",x"06",x"89",x"84",x"60",x"42",x"06",x"60",x"88",x"04",x"40",x"20",x"40",x"84",x"60",x"42",x"06",x"88",x"89",x"85",x"89",x"06",x"20",x"c0",x"38",x"04",x"40",x"40",x"20",x"40",x"84",x"60",x"42",x"06",x"88",x"89",x"85",x"89",x"06",x"20",x"c0",x"38",x"04",x"40",x"40",x"20",x"40",x"84",x"60",x"42",x"06",x"89",x"89",x"06",x"20",x"40",x"05",x"42",x"06",x"88",x"89",x"05",x"60",x"04",x"38",x"10",x"40",x"ff",x"04",x"40",x"0c",x"40",x"40",x"98",x"18",x"30",x"5f",x"90",x"90",x"0c",x"40",x"20",x"40",x"0c",x"60",x"04",x"40",x"40",x"0c",x"40",x"c7",x"38",x"89",x"c6",x"38",x"40",x"40",x"50",x"38",x"10",x"40",x"ff",x"04",x"40",x"0c",x"60",x"04",x"40",x"40",x"98",x"18",x"30",x"70",x"38",x"98",x"04",x"cf",x"38",x"30",x"f5",x"70",x"98",x"04",x"cf",x"38",x"30",x"de",x"10",x"40",x"40",x"40",x"60",x"40",x"60",x"40",x"60",x"40",x"60",x"80",x"0c",x"60",x"40",x"60",x"40",x"60",x"80",x"90",x"50",x"60",x"40",x"38",x"40",x"62",x"41",x"70",x"ff",x"70",x"40",x"05",x"9a",x"80",x"38",x"c1",x"38",x"c0",x"38",x"38",x"0c",x"38",x"c2",x"38",x"c0",x"38",x"38",x"0c",x"38",x"c1",x"38",x"4a",x"70",x"38",x"c0",x"38",x"49",x"80",x"70",x"60",x"47",x"9a",x"8b",x"38",x"00",x"40",x"40",x"04",x"ce",x"38",x"38",x"04",x"c3",x"38",x"60",x"40",x"50",x"80",x"80",x"90",x"18",x"40",x"c0",x"38",x"05",x"82",x"1a",x"62",x"42",x"45",x"80",x"90",x"80",x"90",x"80",x"9a",x"80",x"84",x"70",x"c4",x"38",x"9a",x"8b",x"38",x"00",x"40",x"40",x"04",x"ce",x"38",x"38",x"60",x"40",x"60",x"40",x"60",x"40",x"44",x"7f",x"20",x"c2",x"38",x"60",x"40",x"80",x"50",x"80",x"80",x"90",x"18",x"40",x"80",x"90",x"60",x"45",x"0c",x"05",x"66",x"42",x"41",x"80",x"98",x"9a",x"50",x"60",x"40",x"40",x"0c",x"70",x"c3",x"38",x"c5",x"38",x"ce",x"38",x"c0",x"38",x"40",x"80",x"98",x"74",x"80",x"90",x"47",x"67",x"47",x"66",x"42",x"66",x"42",x"cb",x"38",x"45",x"66",x"42",x"66",x"42",x"c7",x"38",x"60",x"40",x"05",x"60",x"40",x"38",x"ce",x"38",x"c1",x"38",x"c0",x"38",x"40",x"71",x"60",x"40",x"50",x"80",x"80",x"90",x"18",x"60",x"40",x"40",x"40",x"80",x"98",x"ca",x"38",x"80",x"98",x"c1",x"38",x"60",x"40",x"05",x"60",x"40",x"38",x"c0",x"38",x"40",x"80",x"90",x"7f",x"66",x"60",x"40",x"04",x"40",x"60",x"40",x"18",x"60",x"40",x"42",x"c2",x"38",x"60",x"40",x"60",x"40",x"ff",x"04",x"c0",x"38",x"40",x"60",x"40",x"73",x"84",x"89",x"00",x"1a",x"92",x"92",x"92",x"9a",x"89",x"04",x"00",x"92",x"1a",x"40",x"40",x"40",x"40",x"00",x"1a",x"40",x"92",x"92",x"9a",x"89",x"04",x"00",x"92",x"1a",x"40",x"40",x"40",x"40",x"00",x"1a",x"40",x"92",x"92",x"9a",x"89",x"04",x"00",x"92",x"1a",x"40",x"80",x"98",x"04",x"c0",x"38",x"40",x"80",x"98",x"61",x"44",x"c1",x"38",x"0c",x"0c",x"40",x"9a",x"00",x"cf",x"38",x"c0",x"38",x"41",x"8c",x"72",x"40",x"12",x"60",x"40",x"60",x"40",x"1a",x"c1",x"38",x"40",x"00",x"40",x"66",x"49",x"8c",x"76",x"60",x"40",x"20",x"cb",x"38",x"40",x"00",x"12",x"cd",x"38",x"0c",x"40",x"00",x"1a",x"40",x"cb",x"38",x"60",x"40",x"50",x"38",x"c0",x"38",x"38",x"40",x"80",x"90",x"80",x"0c",x"40",x"ff",x"70",x"1a",x"0c",x"40",x"80",x"98",x"0c",x"40",x"ff",x"ff",x"8c",x"04",x"00",x"12",x"60",x"40",x"40",x"60",x"45",x"80",x"98",x"71",x"60",x"42",x"cf",x"38",x"60",x"40",x"60",x"40",x"40",x"c0",x"38",x"40",x"82",x"0c",x"80",x"90",x"0c",x"40",x"80",x"98",x"00",x"60",x"40",x"40",x"67",x"41",x"80",x"98",x"7f",x"04",x"40",x"60",x"40",x"60",x"40",x"6f",x"42",x"70",x"60",x"40",x"05",x"90",x"90",x"c0",x"38",x"60",x"40",x"71",x"40",x"0c",x"40",x"80",x"98",x"71",x"60",x"42",x"cf",x"38",x"60",x"40",x"60",x"40",x"40",x"c0",x"38",x"40",x"0c",x"0c",x"40",x"80",x"98",x"7f",x"04",x"40",x"60",x"40",x"20",x"18",x"c9",x"38",x"c6",x"38",x"60",x"40",x"70",x"04",x"05",x"60",x"40",x"80",x"90",x"80",x"98",x"80",x"80",x"90",x"80",x"98",x"71",x"04",x"c0",x"38",x"40",x"7f",x"60",x"40",x"ca",x"38",x"04",x"ce",x"38",x"60",x"40",x"40",x"80",x"98",x"7f",x"04",x"40",x"60",x"40",x"60",x"41",x"ff",x"1a",x"60",x"42",x"0c",x"60",x"42",x"80",x"9a",x"60",x"42",x"5f",x"60",x"41",x"80",x"98",x"71",x"20",x"60",x"41",x"80",x"98",x"07",x"45",x"c1",x"38",x"72",x"20",x"80",x"90",x"80",x"90",x"cf",x"38",x"60",x"40",x"06",x"80",x"90",x"80",x"98",x"00",x"40",x"72",x"50",x"60",x"40",x"60",x"42",x"40",x"80",x"50",x"40",x"12",x"80",x"c8",x"38",x"ca",x"38",x"50",x"c7",x"38",x"60",x"40",x"60",x"40",x"38",x"60",x"40",x"40",x"80",x"98",x"c6",x"38",x"80",x"98",x"7f",x"40",x"50",x"80",x"80",x"90",x"18",x"80",x"c2",x"38",x"80",x"c0",x"38",x"60",x"40",x"40",x"60",x"40",x"70",x"60",x"40",x"80",x"90",x"80",x"98",x"ca",x"38",x"60",x"41",x"70",x"60",x"40",x"70",x"04",x"60",x"40",x"60",x"40",x"60",x"40",x"40",x"6f",x"c0",x"38",x"80",x"98",x"72",x"05",x"60",x"40",x"04",x"60",x"40",x"1a",x"60",x"40",x"c3",x"38",x"60",x"40",x"70",x"72",x"40",x"80",x"90",x"80",x"98",x"5f",x"40",x"70",x"40",x"60",x"42",x"ca",x"38",x"40",x"8a",x"04",x"20",x"60",x"40",x"40",x"20",x"40",x"5f",x"60",x"40",x"c2",x"38",x"0c",x"60",x"70",x"45",x"9a",x"50",x"92",x"50",x"ce",x"38",x"80",x"98",x"0c",x"c8",x"38",x"20",x"20",x"40",x"5f",x"61",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"40",x"80",x"72",x"40",x"0c",x"40",x"40",x"80",x"90",x"70",x"6f",x"46",x"8c",x"00",x"07",x"12",x"ce",x"38",x"60",x"43",x"70",x"80",x"98",x"0c",x"c7",x"38",x"06",x"20",x"72",x"c9",x"38",x"80",x"98",x"50",x"40",x"80",x"98",x"72",x"70",x"c0",x"38",x"80",x"90",x"70",x"05",x"64",x"c0",x"38",x"40",x"04",x"80",x"90",x"80",x"90",x"80",x"90",x"66",x"42",x"0c",x"40",x"80",x"90",x"cf",x"38",x"60",x"40",x"ce",x"38",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"60",x"40",x"60",x"40",x"ce",x"38",x"40",x"6f",x"45",x"07",x"46",x"80",x"8c",x"80",x"90",x"80",x"8c",x"90",x"8c",x"90",x"80",x"90",x"80",x"98",x"80",x"98",x"c9",x"38",x"40",x"c0",x"38",x"60",x"41",x"72",x"60",x"40",x"60",x"40",x"60",x"80",x"98",x"c0",x"38",x"38",x"80",x"92",x"40",x"80",x"60",x"42",x"80",x"98",x"0c",x"50",x"50",x"50",x"cf",x"38",x"60",x"41",x"76",x"20",x"60",x"40",x"98",x"60",x"41",x"80",x"98",x"80",x"98",x"70",x"cf",x"38",x"60",x"41",x"70",x"38",x"40",x"80",x"6f",x"60",x"40",x"43",x"80",x"98",x"72",x"20",x"12",x"38",x"60",x"40",x"00",x"0c",x"c1",x"38",x"60",x"40",x"70",x"40",x"c0",x"38",x"cf",x"38",x"76",x"40",x"60",x"40",x"0c",x"40",x"70",x"40",x"53",x"40",x"40",x"70",x"12",x"60",x"40",x"60",x"40",x"80",x"98",x"60",x"42",x"60",x"60",x"40",x"41",x"40",x"50",x"64",x"47",x"60",x"42",x"62",x"42",x"4e",x"f0",x"64",x"42",x"66",x"41",x"0c",x"40",x"40",x"c0",x"38",x"0c",x"ce",x"38",x"20",x"c1",x"38",x"20",x"60",x"92",x"ce",x"38",x"38",x"40",x"12",x"20",x"ca",x"38",x"ca",x"38",x"80",x"0c",x"1a",x"60",x"41",x"70",x"50",x"c0",x"38",x"60",x"41",x"70",x"c6",x"38",x"38",x"50",x"60",x"42",x"64",x"42",x"66",x"41",x"0c",x"9a",x"80",x"63",x"42",x"62",x"41",x"80",x"07",x"42",x"00",x"60",x"82",x"80",x"80",x"70",x"40",x"80",x"9a",x"80",x"98",x"80",x"98",x"80",x"0c",x"40",x"60",x"c1",x"38",x"40",x"40",x"c0",x"38",x"0c",x"ce",x"38",x"20",x"82",x"04",x"c4",x"38",x"c0",x"38",x"38",x"60",x"80",x"98",x"00",x"20",x"0c",x"c2",x"38",x"60",x"40",x"7f",x"60",x"40",x"38",x"80",x"98",x"ff",x"04",x"c1",x"38",x"60",x"40",x"50",x"60",x"40",x"04",x"c4",x"38",x"c0",x"38",x"38",x"60",x"40",x"60",x"40",x"40",x"04",x"ca",x"38",x"7f",x"60",x"40",x"38",x"80",x"98",x"80",x"98",x"70",x"c1",x"38",x"60",x"40",x"38",x"80",x"0c",x"50",x"1a",x"c0",x"38",x"38",x"60",x"40",x"0c",x"c2",x"38",x"72",x"c3",x"38",x"80",x"c1",x"38",x"20",x"40",x"40",x"90",x"8c",x"90",x"80",x"98",x"80",x"98",x"c7",x"38",x"40",x"c0",x"38",x"60",x"41",x"72",x"60",x"40",x"60",x"40",x"60",x"42",x"43",x"73",x"12",x"44",x"cb",x"38",x"73",x"92",x"80",x"c9",x"38",x"20",x"40",x"40",x"98",x"70",x"c6",x"38",x"73",x"70",x"40",x"50",x"c0",x"38",x"38",x"50",x"98",x"82",x"07",x"45",x"1a",x"c2",x"38",x"80",x"50",x"40",x"60",x"42",x"4e",x"98",x"50",x"07",x"41",x"72",x"50",x"12",x"9a",x"60",x"42",x"4d",x"50",x"40",x"70",x"80",x"9a",x"60",x"42",x"80",x"0c",x"40",x"18",x"40",x"60",x"41",x"38",x"10",x"40",x"40",x"60",x"41",x"98",x"98",x"98",x"18",x"40",x"38",x"58",x"90",x"90",x"90",x"0c",x"71",x"40",x"04",x"c0",x"38",x"84",x"74",x"40",x"60",x"42",x"f1",x"70",x"40",x"c6",x"38",x"70",x"60",x"42",x"6f",x"43",x"41",x"70",x"60",x"42",x"5f",x"42",x"70",x"72",x"20",x"38",x"40",x"8a",x"04",x"04",x"40",x"20",x"90",x"84",x"60",x"40",x"41",x"41",x"60",x"42",x"41",x"5f",x"40",x"38",x"40",x"38",x"40",x"c0",x"38",x"0c",x"40",x"90",x"90",x"60",x"05",x"40",x"42",x"70",x"90",x"8c",x"0c",x"00",x"40",x"c2",x"38",x"40",x"1a",x"40",x"0c",x"ce",x"38",x"50",x"cc",x"38",x"38",x"70",x"92",x"90",x"0c",x"40",x"c0",x"38",x"90",x"98",x"98",x"98",x"82",x"71",x"60",x"41",x"60",x"44",x"41",x"0c",x"0c",x"40",x"00",x"40",x"5f",x"40",x"40",x"60",x"42",x"12",x"98",x"0c",x"c2",x"38",x"c0",x"38",x"38",x"92",x"73",x"50",x"38",x"c0",x"38",x"12",x"98",x"98",x"71",x"60",x"41",x"60",x"44",x"42",x"98",x"ff",x"0c",x"04",x"c6",x"38",x"7f",x"38",x"98",x"07",x"44",x"0c",x"20",x"0c",x"0c",x"40",x"0c",x"40",x"0c",x"c1",x"38",x"0c",x"8c",x"60",x"1a",x"50",x"43",x"00",x"c0",x"38",x"38",x"72",x"0c",x"40",x"80",x"40",x"0c",x"40",x"40",x"40",x"57",x"38",x"70",x"90",x"90",x"f6",x"90",x"98",x"90",x"40",x"98",x"18",x"30",x"5c",x"90",x"90",x"90",x"90",x"0c",x"70",x"40",x"40",x"40",x"70",x"c0",x"38",x"98",x"98",x"70",x"c2",x"38",x"70",x"43",x"70",x"40",x"70",x"c0",x"38",x"70",x"84",x"98",x"74",x"43",x"0c",x"40",x"40",x"10",x"41",x"70",x"80",x"70",x"98",x"8c",x"c9",x"38",x"40",x"40",x"70",x"98",x"90",x"98",x"90",x"c1",x"38",x"cd",x"38",x"40",x"80",x"90",x"98",x"98",x"90",x"a4",x"70",x"ce",x"38",x"40",x"c3",x"38",x"9e",x"75",x"70",x"90",x"90",x"ce",x"38",x"a4",x"70",x"c5",x"38",x"c6",x"38",x"70",x"92",x"98",x"90",x"98",x"90",x"c8",x"38",x"40",x"40",x"98",x"5f",x"c7",x"38",x"40",x"c0",x"38",x"40",x"98",x"0c",x"50",x"50",x"cf",x"38",x"40",x"40",x"40",x"98",x"98",x"70",x"ca",x"38",x"70",x"41",x"70",x"40",x"70",x"40",x"40",x"40",x"60",x"c0",x"38",x"98",x"05",x"04",x"c0",x"38",x"38",x"40",x"40",x"60",x"70",x"40",x"40",x"40",x"40",x"0c",x"60",x"70",x"40",x"ca",x"38",x"40",x"98",x"0c",x"40",x"45",x"90",x"98",x"90",x"98",x"98",x"0c",x"38",x"40",x"40",x"38",x"40",x"40",x"98",x"0c",x"98",x"90",x"10",x"c0",x"38",x"98",x"00",x"ca",x"38",x"20",x"40",x"90",x"c6",x"38",x"40",x"07",x"40",x"48",x"98",x"0c",x"60",x"70",x"ca",x"38",x"40",x"c5",x"38",x"40",x"98",x"98",x"ca",x"38",x"40",x"0c",x"50",x"c0",x"38",x"40",x"ca",x"38",x"40",x"c0",x"38",x"38",x"98",x"73",x"0c",x"50",x"98",x"42",x"70",x"45",x"98",x"70",x"40",x"38",x"40",x"92",x"5f",x"38",x"c3",x"38",x"07",x"4a",x"4d",x"12",x"18",x"10",x"41",x"07",x"4a",x"12",x"4c",x"70",x"98",x"98",x"98",x"18",x"30",x"00",x"70",x"90",x"90",x"98",x"90",x"98",x"90",x"c1",x"38",x"40",x"51",x"38",x"5e",x"40",x"90",x"90",x"90",x"98",x"90",x"ce",x"38",x"40",x"51",x"38",x"5e",x"40",x"90",x"90",x"90",x"98",x"90",x"cb",x"38",x"40",x"51",x"38",x"38",x"38",x"38",x"30",x"00",x"10",x"40",x"40",x"0c",x"60",x"70",x"40",x"98",x"18",x"30",x"00",x"12",x"38",x"12",x"38",x"84",x"60",x"41",x"42",x"0c",x"c7",x"38",x"50",x"84",x"60",x"41",x"40",x"0c",x"c4",x"38",x"40",x"04",x"40",x"88",x"05",x"4a",x"10",x"40",x"40",x"40",x"51",x"ce",x"38",x"38",x"50",x"60",x"47",x"60",x"42",x"12",x"50",x"cf",x"38",x"38",x"89",x"ff",x"10",x"40",x"fc",x"00",x"c4",x"38",x"c0",x"38",x"40",x"8f",x"7f",x"20",x"20",x"60",x"41",x"45",x"7f",x"06",x"10",x"40",x"43",x"63",x"44",x"fb",x"00",x"89",x"84",x"60",x"42",x"06",x"84",x"90",x"0c",x"40",x"0c",x"38",x"90",x"80",x"70",x"70",x"38",x"70",x"04",x"90",x"98",x"18",x"50",x"38",x"10",x"40",x"40",x"7f",x"ff",x"7f",x"40",x"20",x"20",x"20",x"ef",x"6f",x"c0",x"38",x"6f",x"c0",x"38",x"c0",x"38",x"84",x"84",x"60",x"41",x"7f",x"20",x"20",x"ef",x"6f",x"c0",x"38",x"6f",x"c0",x"38",x"c0",x"38",x"04",x"c0",x"38",x"70",x"c0",x"38",x"70",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c1",x"38",x"60",x"0c",x"0c",x"40",x"70",x"60",x"42",x"70",x"f0",x"60",x"49",x"70",x"42",x"0c",x"60",x"41",x"88",x"70",x"05",x"ce",x"38",x"60",x"86",x"05",x"c3",x"38",x"20",x"70",x"86",x"06",x"f8",x"70",x"c0",x"38",x"70",x"42",x"0c",x"ca",x"38",x"05",x"c0",x"38",x"0c",x"c8",x"38",x"20",x"c0",x"38",x"40",x"85",x"0c",x"0c",x"42",x"70",x"07",x"47",x"70",x"c0",x"38",x"c0",x"38",x"0c",x"c0",x"38",x"c0",x"38",x"0c",x"41",x"0c",x"41",x"0c",x"40",x"40",x"84",x"8f",x"7f",x"84",x"c0",x"38",x"40",x"40",x"90",x"60",x"42",x"89",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"89",x"46",x"89",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"72",x"40",x"20",x"40",x"0c",x"40",x"0c",x"0c",x"20",x"40",x"40",x"40",x"20",x"60",x"60",x"c1",x"38",x"40",x"40",x"40",x"90",x"60",x"42",x"89",x"90",x"0c",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"40",x"38",x"40",x"90",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"72",x"40",x"20",x"40",x"c0",x"38",x"0c",x"82",x"88",x"89",x"88",x"07",x"80",x"70",x"20",x"41",x"0c",x"45",x"82",x"70",x"63",x"47",x"0c",x"90",x"90",x"ca",x"38",x"40",x"74",x"40",x"20",x"c9",x"38",x"20",x"60",x"41",x"70",x"40",x"40",x"98",x"98",x"86",x"80",x"70",x"04",x"40",x"40",x"40",x"40",x"40",x"88",x"80",x"70",x"c0",x"38",x"38",x"20",x"20",x"60",x"04",x"c5",x"38",x"40",x"40",x"70",x"40",x"05",x"85",x"c3",x"38",x"0c",x"70",x"06",x"20",x"03",x"cd",x"38",x"60",x"c1",x"38",x"40",x"c8",x"38",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"40",x"40",x"85",x"0c",x"0c",x"41",x"84",x"84",x"0c",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"72",x"40",x"80",x"0c",x"0c",x"40",x"98",x"0c",x"82",x"ef",x"c1",x"38",x"40",x"60",x"70",x"05",x"40",x"60",x"43",x"70",x"82",x"82",x"0c",x"40",x"c8",x"38",x"60",x"41",x"70",x"40",x"0c",x"40",x"0c",x"20",x"89",x"8f",x"7f",x"40",x"70",x"88",x"05",x"05",x"40",x"88",x"05",x"04",x"c0",x"38",x"0e",x"20",x"c0",x"38",x"70",x"0e",x"0c",x"40",x"40",x"40",x"52",x"38",x"04",x"c1",x"38",x"40",x"88",x"70",x"38",x"c1",x"38",x"88",x"82",x"89",x"88",x"70",x"05",x"30",x"00",x"70",x"10",x"c0",x"38",x"ff",x"7f",x"84",x"f0",x"60",x"47",x"70",x"42",x"0c",x"60",x"41",x"04",x"70",x"c0",x"38",x"70",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c8",x"38",x"20",x"20",x"70",x"c7",x"38",x"20",x"c2",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c2",x"38",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c0",x"38",x"04",x"60",x"41",x"70",x"06",x"60",x"41",x"70",x"0c",x"30",x"00",x"70",x"10",x"c0",x"38",x"ff",x"7f",x"84",x"f0",x"60",x"47",x"70",x"42",x"0c",x"7f",x"cb",x"38",x"70",x"60",x"41",x"70",x"f0",x"60",x"47",x"70",x"42",x"0c",x"60",x"41",x"85",x"85",x"05",x"60",x"42",x"84",x"60",x"45",x"70",x"07",x"49",x"70",x"07",x"45",x"70",x"42",x"42",x"70",x"07",x"47",x"70",x"07",x"43",x"70",x"42",x"0c",x"60",x"c1",x"38",x"06",x"05",x"c0",x"38",x"18",x"50",x"38",x"ff",x"7f",x"70",x"04",x"c0",x"38",x"f0",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c2",x"38",x"60",x"70",x"04",x"c0",x"38",x"f0",x"60",x"47",x"70",x"42",x"0c",x"50",x"38",x"5f",x"70",x"60",x"41",x"70",x"60",x"70",x"20",x"60",x"c0",x"38",x"c0",x"38",x"04",x"cb",x"38",x"70",x"60",x"41",x"70",x"f0",x"60",x"47",x"70",x"42",x"0c",x"60",x"41",x"85",x"85",x"05",x"60",x"42",x"84",x"60",x"45",x"70",x"07",x"49",x"70",x"07",x"45",x"70",x"42",x"42",x"70",x"07",x"47",x"70",x"07",x"43",x"70",x"42",x"0c",x"7f",x"c1",x"38",x"06",x"05",x"c0",x"38",x"18",x"50",x"38",x"5f",x"70",x"60",x"41",x"70",x"60",x"70",x"20",x"60",x"c0",x"38",x"c0",x"38",x"04",x"cb",x"38",x"70",x"60",x"41",x"70",x"f0",x"60",x"47",x"70",x"42",x"0c",x"60",x"41",x"85",x"85",x"05",x"60",x"42",x"84",x"60",x"45",x"70",x"07",x"49",x"70",x"07",x"45",x"70",x"42",x"42",x"70",x"07",x"47",x"70",x"07",x"43",x"70",x"42",x"0c",x"7f",x"c1",x"38",x"06",x"05",x"c0",x"38",x"18",x"50",x"38",x"5f",x"70",x"60",x"41",x"70",x"60",x"70",x"20",x"60",x"c0",x"38",x"c0",x"38",x"04",x"cb",x"38",x"70",x"60",x"41",x"70",x"f0",x"60",x"47",x"70",x"42",x"0c",x"60",x"41",x"85",x"85",x"05",x"60",x"42",x"84",x"60",x"45",x"70",x"07",x"49",x"70",x"07",x"45",x"70",x"42",x"42",x"70",x"07",x"47",x"70",x"07",x"43",x"70",x"42",x"0c",x"7f",x"c1",x"38",x"06",x"05",x"c0",x"38",x"18",x"50",x"38",x"5f",x"70",x"60",x"41",x"70",x"60",x"70",x"20",x"60",x"c0",x"38",x"c0",x"38",x"04",x"60",x"41",x"04",x"70",x"c0",x"38",x"70",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c8",x"38",x"20",x"20",x"70",x"c7",x"38",x"20",x"c2",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c2",x"38",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c0",x"38",x"04",x"7f",x"41",x"70",x"06",x"60",x"41",x"70",x"0c",x"30",x"00",x"0c",x"20",x"70",x"10",x"40",x"40",x"40",x"89",x"90",x"ff",x"04",x"40",x"40",x"8f",x"7f",x"20",x"90",x"90",x"80",x"ef",x"c1",x"38",x"40",x"ef",x"c0",x"38",x"40",x"ff",x"7f",x"40",x"70",x"84",x"c0",x"38",x"70",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c1",x"38",x"60",x"85",x"c0",x"38",x"20",x"70",x"c0",x"38",x"70",x"60",x"c0",x"38",x"98",x"c0",x"38",x"04",x"c2",x"38",x"60",x"0c",x"20",x"40",x"70",x"40",x"40",x"60",x"90",x"89",x"70",x"90",x"88",x"85",x"84",x"73",x"20",x"0c",x"40",x"c8",x"38",x"70",x"82",x"70",x"40",x"89",x"88",x"70",x"85",x"70",x"c5",x"38",x"70",x"82",x"70",x"40",x"89",x"88",x"70",x"85",x"70",x"c2",x"38",x"70",x"82",x"70",x"40",x"89",x"88",x"70",x"80",x"98",x"0c",x"40",x"cf",x"38",x"40",x"70",x"70",x"40",x"8e",x"70",x"0c",x"70",x"70",x"70",x"40",x"90",x"70",x"70",x"cb",x"38",x"40",x"7f",x"01",x"0e",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"c0",x"70",x"20",x"70",x"40",x"90",x"70",x"70",x"40",x"40",x"98",x"88",x"70",x"20",x"81",x"98",x"70",x"40",x"0e",x"70",x"90",x"7f",x"40",x"20",x"c2",x"38",x"40",x"70",x"20",x"81",x"70",x"20",x"40",x"20",x"40",x"40",x"60",x"82",x"98",x"80",x"c5",x"38",x"40",x"0c",x"40",x"40",x"40",x"98",x"70",x"0f",x"40",x"45",x"f0",x"70",x"20",x"60",x"41",x"06",x"60",x"41",x"c8",x"38",x"40",x"40",x"40",x"0c",x"40",x"40",x"40",x"40",x"98",x"70",x"88",x"03",x"40",x"60",x"ef",x"c0",x"38",x"40",x"98",x"60",x"43",x"46",x"98",x"0e",x"81",x"70",x"70",x"47",x"70",x"c0",x"38",x"c0",x"38",x"8f",x"7f",x"40",x"05",x"40",x"01",x"85",x"05",x"40",x"06",x"60",x"41",x"70",x"40",x"70",x"40",x"98",x"85",x"60",x"41",x"c9",x"38",x"20",x"c7",x"38",x"8f",x"6f",x"47",x"60",x"42",x"89",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"89",x"ca",x"38",x"60",x"70",x"41",x"85",x"60",x"42",x"70",x"38",x"60",x"70",x"40",x"40",x"40",x"0c",x"53",x"38",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"89",x"85",x"80",x"0c",x"cf",x"38",x"70",x"82",x"98",x"8f",x"6f",x"4a",x"47",x"90",x"60",x"42",x"89",x"90",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"89",x"47",x"90",x"90",x"90",x"c1",x"38",x"40",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"89",x"85",x"80",x"0c",x"cd",x"38",x"80",x"0c",x"90",x"c9",x"38",x"10",x"40",x"40",x"0c",x"40",x"20",x"20",x"40",x"20",x"20",x"40",x"86",x"98",x"98",x"18",x"40",x"82",x"50",x"38",x"10",x"40",x"7f",x"c0",x"38",x"8f",x"7f",x"60",x"04",x"40",x"ff",x"04",x"70",x"63",x"47",x"73",x"20",x"40",x"41",x"70",x"c1",x"38",x"40",x"40",x"0c",x"40",x"0c",x"40",x"0c",x"30",x"00",x"40",x"40",x"70",x"70",x"60",x"45",x"60",x"45",x"89",x"88",x"f1",x"05",x"70",x"82",x"05",x"20",x"30",x"00",x"0c",x"70",x"90",x"60",x"42",x"89",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"71",x"40",x"20",x"82",x"70",x"40",x"90",x"70",x"06",x"40",x"f0",x"50",x"40",x"0c",x"30",x"00",x"04",x"c1",x"38",x"40",x"20",x"41",x"60",x"42",x"72",x"20",x"20",x"20",x"20",x"70",x"0c",x"38",x"10",x"40",x"40",x"0c",x"40",x"8b",x"98",x"82",x"98",x"18",x"30",x"00",x"10",x"40",x"40",x"40",x"86",x"80",x"70",x"04",x"40",x"40",x"40",x"90",x"89",x"04",x"60",x"84",x"04",x"40",x"40",x"40",x"40",x"40",x"47",x"98",x"5f",x"40",x"48",x"c9",x"38",x"60",x"70",x"60",x"20",x"42",x"70",x"f0",x"60",x"49",x"70",x"42",x"0c",x"60",x"41",x"88",x"70",x"20",x"40",x"84",x"70",x"60",x"42",x"70",x"f0",x"60",x"49",x"70",x"42",x"0c",x"60",x"41",x"88",x"70",x"05",x"40",x"70",x"40",x"40",x"70",x"90",x"0c",x"cf",x"38",x"40",x"40",x"40",x"98",x"88",x"85",x"98",x"90",x"70",x"20",x"0c",x"40",x"40",x"90",x"80",x"70",x"98",x"85",x"f0",x"04",x"20",x"0c",x"90",x"70",x"40",x"40",x"90",x"0e",x"70",x"40",x"0c",x"40",x"98",x"c7",x"38",x"40",x"40",x"0e",x"0e",x"40",x"70",x"20",x"40",x"20",x"60",x"84",x"98",x"60",x"98",x"98",x"00",x"40",x"d0",x"c3",x"38",x"43",x"f0",x"70",x"20",x"60",x"41",x"98",x"85",x"60",x"41",x"47",x"8e",x"89",x"85",x"01",x"01",x"40",x"ef",x"c0",x"38",x"38",x"c0",x"38",x"38",x"40",x"60",x"88",x"04",x"c8",x"38",x"40",x"05",x"c5",x"38",x"20",x"c1",x"38",x"60",x"70",x"cb",x"38",x"60",x"70",x"40",x"70",x"40",x"40",x"20",x"64",x"40",x"49",x"70",x"40",x"98",x"85",x"60",x"41",x"c6",x"38",x"20",x"c0",x"38",x"40",x"70",x"60",x"cf",x"38",x"c6",x"38",x"40",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"40",x"40",x"0c",x"0c",x"c0",x"38",x"90",x"0c",x"40",x"20",x"90",x"cf",x"38",x"60",x"41",x"70",x"40",x"40",x"40",x"40",x"0c",x"40",x"98",x"0c",x"90",x"98",x"98",x"05",x"0c",x"40",x"ca",x"38",x"40",x"70",x"70",x"70",x"c0",x"38",x"98",x"60",x"41",x"70",x"42",x"0c",x"40",x"70",x"8e",x"81",x"80",x"70",x"05",x"c1",x"38",x"70",x"0e",x"40",x"70",x"38",x"0c",x"40",x"40",x"40",x"0c",x"30",x"89",x"90",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"72",x"40",x"20",x"40",x"0c",x"40",x"98",x"0c",x"0c",x"20",x"60",x"c0",x"38",x"38",x"40",x"c7",x"38",x"40",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"40",x"38",x"40",x"40",x"40",x"89",x"90",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"72",x"40",x"20",x"40",x"0c",x"40",x"90",x"80",x"0c",x"20",x"40",x"40",x"00",x"89",x"89",x"8b",x"10",x"20",x"80",x"7f",x"20",x"20",x"8b",x"8b",x"89",x"00",x"20",x"20",x"20",x"20",x"00",x"40",x"05",x"40",x"40",x"0c",x"50",x"38",x"80",x"70",x"90",x"06",x"40",x"98",x"18",x"30",x"00",x"60",x"42",x"60",x"42",x"89",x"05",x"40",x"89",x"05",x"40",x"89",x"85",x"89",x"05",x"40",x"89",x"05",x"86",x"d5",x"75",x"40",x"82",x"89",x"05",x"40",x"b3",x"73",x"84",x"89",x"04",x"40",x"00",x"20",x"40",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"81",x"70",x"20",x"20",x"40",x"40",x"20",x"c6",x"38",x"41",x"30",x"71",x"82",x"50",x"88",x"c3",x"38",x"20",x"80",x"70",x"40",x"40",x"40",x"60",x"05",x"20",x"40",x"20",x"20",x"20",x"41",x"88",x"85",x"0c",x"38",x"10",x"40",x"40",x"0c",x"40",x"8b",x"98",x"82",x"98",x"18",x"30",x"00",x"33",x"e7",x"be",x"56",x"07",x"39",x"8e",x"00",x"62",x"62",x"62",x"62",x"62",x"62",x"62",x"62",x"62",x"62",x"62",x"62",x"62",x"62",x"62",x"62",x"61",x"00",x"70",x"61",x"36",x"65",x"72",x"63",x"75",x"61",x"65",x"73",x"72",x"72",x"72",x"00",x"76",x"64",x"6f",x"75",x"61",x"65",x"73",x"72",x"72",x"72",x"00",x"66",x"20",x"65",x"69",x"72",x"70",x"6d",x"72",x"6f",x"6f",x"61",x"0a",x"20",x"66",x"61",x"20",x"20",x"61",x"65",x"66",x"63",x"6d",x"2e",x"4b",x"6c",x"74",x"20",x"20",x"61",x"65",x"66",x"63",x"6d",x"2e",x"25",x"52",x"21",x"73",x"72",x"78",x"78",x"73",x"6c",x"65",x"25",x"0a",x"75",x"52",x"20",x"72",x"63",x"30",x"34",x"20",x"75",x"62",x"78",x"78",x"25",x"52",x"21",x"61",x"63",x"30",x"34",x"20",x"75",x"62",x"78",x"78",x"6f",x"61",x"53",x"20",x"3a",x"75",x"6f",x"20",x"6b",x"20",x"3a",x"75",x"6f",x"20",x"65",x"65",x"3a",x"0a",x"65",x"69",x"2f",x"20",x"20",x"00",x"4f",x"4d",x"20",x"63",x"20",x"20",x"6c",x"74",x"20",x"73",x"72",x"76",x"64",x"73",x"21",x"74",x"74",x"73",x"20",x"3a",x"75",x"6f",x"6c",x"76",x"69",x"3a",x"0a",x"43",x"2e",x"6f",x"74",x"65",x"61",x"33",x"28",x"73",x"4c",x"45",x"2f",x"61",x"43",x"69",x"20",x"67",x"20",x"73",x"65",x"79",x"63",x"6f",x"3a",x"0a",x"41",x"73",x"63",x"20",x"20",x"20",x"78",x"78",x"25",x"72",x"73",x"20",x"20",x"78",x"78",x"25",x"72",x"74",x"20",x"20",x"78",x"78",x"25",x"72",x"61",x"20",x"20",x"78",x"78",x"25",x"72",x"6e",x"20",x"20",x"78",x"78",x"6f",x"63",x"70",x"74",x"20",x"69",x"65",x"53",x"72",x"6d",x"78",x"6f",x"75",x"6e",x"65",x"74",x"20",x"65",x"00",x"65",x"6b",x"30",x"25",x"20",x"25",x"2f",x"00",x"6f",x"64",x"63",x"0a",x"6e",x"20",x"69",x"65",x"65",x"69",x"66",x"74",x"65",x"65",x"61",x"73",x"6c",x"65",x"6d",x"65",x"74",x"65",x"74",x"6e",x"6b",x"6e",x"61",x"72",x"00",x"33",x"46",x"2e",x"54",x"54",x"65",x"33",x"65",x"00",x"30",x"33",x"31",x"2d",x"38",x"38",x"2b",x"65",x"00",x"35",x"30",x"32",x"30",x"31",x"37",x"2b",x"34",x"00",x"32",x"33",x"38",x"2b",x"00",x"4c",x"30",x"34",x"38",x"63",x"67",x"6b",x"6f",x"73",x"77",x"00",x"33",x"37",x"42",x"46",x"4a",x"4e",x"52",x"56",x"5a",x"00",x"5e",x"5e",x"5e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
 shared variable RAM2: RAM_TABLE := RAM_TABLE'(
x"00",x"01",x"be",x"f2",x"95",x"21",x"41",x"02",x"00",x"01",x"04",x"cf",x"00",x"41",x"11",x"00",x"02",x"04",x"14",x"53",x"20",x"43",x"00",x"00",x"00",x"0a",x"41",x"12",x"02",x"ff",x"11",x"10",x"01",x"10",x"10",x"0f",x"4f",x"5f",x"6f",x"1f",x"26",x"13",x"00",x"01",x"00",x"f1",x"20",x"10",x"03",x"21",x"04",x"71",x"01",x"00",x"20",x"3f",x"22",x"14",x"18",x"02",x"96",x"9f",x"29",x"00",x"29",x"84",x"9f",x"0d",x"10",x"16",x"65",x"01",x"00",x"46",x"40",x"11",x"00",x"e0",x"3f",x"61",x"36",x"4d",x"10",x"16",x"65",x"01",x"00",x"46",x"c0",x"65",x"3f",x"34",x"ff",x"f1",x"0d",x"10",x"ff",x"01",x"00",x"18",x"f1",x"12",x"3f",x"23",x"0c",x"10",x"14",x"0f",x"10",x"0f",x"4f",x"34",x"08",x"6f",x"42",x"fe",x"16",x"42",x"fe",x"16",x"6f",x"5f",x"4f",x"df",x"d0",x"03",x"00",x"31",x"ff",x"03",x"08",x"08",x"00",x"98",x"82",x"83",x"08",x"73",x"11",x"22",x"11",x"21",x"d0",x"32",x"22",x"21",x"d0",x"0f",x"4f",x"5f",x"6f",x"1f",x"51",x"11",x"18",x"18",x"10",x"00",x"00",x"10",x"00",x"0a",x"00",x"1e",x"00",x"26",x"14",x"1f",x"01",x"1c",x"62",x"60",x"10",x"10",x"04",x"02",x"02",x"60",x"10",x"10",x"09",x"80",x"10",x"10",x"02",x"94",x"99",x"29",x"00",x"80",x"44",x"04",x"ff",x"a0",x"49",x"10",x"02",x"20",x"10",x"54",x"42",x"20",x"10",x"09",x"00",x"25",x"22",x"22",x"10",x"29",x"10",x"10",x"04",x"22",x"04",x"40",x"10",x"10",x"09",x"b4",x"2f",x"29",x"02",x"00",x"42",x"95",x"25",x"00",x"1a",x"22",x"e2",x"a2",x"20",x"10",x"14",x"00",x"2f",x"2f",x"e0",x"03",x"07",x"3f",x"11",x"12",x"04",x"00",x"3f",x"51",x"01",x"01",x"15",x"10",x"15",x"21",x"7f",x"37",x"31",x"27",x"21",x"21",x"07",x"60",x"10",x"10",x"20",x"10",x"00",x"61",x"26",x"22",x"12",x"00",x"66",x"80",x"10",x"10",x"14",x"e0",x"10",x"16",x"11",x"21",x"00",x"66",x"80",x"10",x"06",x"00",x"ff",x"f1",x"02",x"04",x"11",x"1e",x"66",x"06",x"ff",x"7f",x"15",x"04",x"04",x"04",x"04",x"21",x"71",x"42",x"cd",x"10",x"65",x"60",x"10",x"00",x"14",x"15",x"11",x"4d",x"10",x"14",x"e0",x"10",x"00",x"6f",x"5f",x"41",x"0c",x"0f",x"10",x"12",x"17",x"f7",x"00",x"40",x"03",x"00",x"ff",x"f2",x"73",x"77",x"27",x"00",x"e0",x"33",x"40",x"10",x"10",x"40",x"10",x"22",x"04",x"01",x"60",x"10",x"10",x"03",x"ff",x"d0",x"31",x"10",x"d0",x"03",x"60",x"10",x"10",x"12",x"23",x"20",x"10",x"d0",x"02",x"d0",x"4f",x"11",x"4f",x"5f",x"6f",x"3f",x"2f",x"1f",x"09",x"00",x"00",x"10",x"08",x"02",x"0a",x"1f",x"01",x"20",x"28",x"8f",x"07",x"00",x"10",x"00",x"29",x"3f",x"0a",x"00",x"18",x"00",x"0b",x"00",x"0a",x"00",x"1b",x"0a",x"b3",x"10",x"a0",x"10",x"80",x"10",x"fa",x"93",x"14",x"60",x"10",x"10",x"e0",x"2f",x"0b",x"00",x"12",x"0a",x"24",x"20",x"18",x"ff",x"80",x"af",x"86",x"b4",x"04",x"04",x"18",x"1c",x"10",x"40",x"10",x"10",x"41",x"68",x"c0",x"14",x"10",x"52",x"f8",x"ff",x"3f",x"00",x"10",x"28",x"14",x"02",x"12",x"60",x"10",x"10",x"20",x"60",x"10",x"28",x"10",x"28",x"1f",x"2a",x"20",x"fe",x"1f",x"12",x"1f",x"11",x"1f",x"1f",x"19",x"fe",x"6f",x"5f",x"4f",x"df",x"d0",x"ed",x"10",x"31",x"72",x"71",x"32",x"31",x"31",x"02",x"10",x"04",x"04",x"04",x"04",x"31",x"d0",x"00",x"df",x"0c",x"42",x"08",x"04",x"14",x"54",x"19",x"03",x"48",x"39",x"03",x"01",x"04",x"04",x"02",x"00",x"31",x"02",x"05",x"00",x"7b",x"9f",x"5b",x"00",x"94",x"10",x"94",x"84",x"7f",x"0c",x"02",x"00",x"87",x"3f",x"83",x"e8",x"10",x"9f",x"00",x"10",x"14",x"00",x"0a",x"8b",x"1b",x"00",x"7e",x"5e",x"00",x"52",x"83",x"06",x"05",x"03",x"63",x"53",x"53",x"34",x"38",x"7f",x"78",x"b8",x"37",x"e7",x"10",x"2a",x"ff",x"64",x"02",x"00",x"3f",x"1f",x"ff",x"f2",x"05",x"4d",x"10",x"02",x"f3",x"78",x"17",x"00",x"89",x"57",x"37",x"96",x"79",x"66",x"07",x"40",x"10",x"42",x"03",x"fc",x"6f",x"5f",x"4f",x"df",x"d0",x"8f",x"04",x"0c",x"83",x"08",x"80",x"10",x"af",x"4b",x"80",x"10",x"87",x"38",x"14",x"04",x"41",x"18",x"32",x"22",x"21",x"4f",x"71",x"d0",x"0f",x"4f",x"14",x"08",x"04",x"54",x"64",x"64",x"64",x"64",x"05",x"00",x"41",x"0d",x"10",x"38",x"18",x"14",x"41",x"8d",x"10",x"38",x"18",x"14",x"06",x"00",x"14",x"16",x"c0",x"10",x"04",x"08",x"0c",x"01",x"d0",x"00",x"f7",x"4f",x"5f",x"6f",x"1f",x"f1",x"23",x"28",x"00",x"48",x"08",x"1f",x"cd",x"10",x"8d",x"10",x"30",x"cd",x"10",x"32",x"0d",x"10",x"34",x"4d",x"10",x"4c",x"8d",x"10",x"01",x"00",x"13",x"50",x"30",x"60",x"10",x"10",x"32",x"01",x"00",x"2f",x"01",x"20",x"10",x"34",x"56",x"1f",x"1f",x"2f",x"80",x"06",x"00",x"1f",x"06",x"e0",x"10",x"34",x"20",x"10",x"61",x"30",x"32",x"34",x"32",x"74",x"08",x"2f",x"2f",x"6f",x"1f",x"11",x"13",x"21",x"31",x"00",x"50",x"01",x"70",x"50",x"00",x"4c",x"02",x"00",x"44",x"21",x"00",x"12",x"07",x"50",x"08",x"3f",x"58",x"48",x"80",x"10",x"3f",x"08",x"2f",x"02",x"00",x"02",x"02",x"12",x"2f",x"08",x"7f",x"08",x"2f",x"02",x"00",x"ff",x"f2",x"12",x"32",x"44",x"60",x"10",x"3c",x"ad",x"10",x"54",x"50",x"71",x"20",x"10",x"32",x"30",x"10",x"21",x"08",x"1f",x"2f",x"14",x"1f",x"0d",x"10",x"50",x"71",x"60",x"10",x"30",x"44",x"1f",x"6d",x"10",x"4c",x"e0",x"10",x"1f",x"a1",x"10",x"4c",x"12",x"1f",x"cd",x"10",x"30",x"fc",x"0d",x"10",x"30",x"0d",x"10",x"00",x"03",x"08",x"1f",x"62",x"3b",x"15",x"40",x"10",x"08",x"1f",x"62",x"7f",x"04",x"3a",x"f1",x"40",x"10",x"51",x"21",x"80",x"10",x"ff",x"08",x"1f",x"62",x"47",x"12",x"40",x"10",x"a1",x"4f",x"2f",x"11",x"01",x"4c",x"30",x"f1",x"08",x"1f",x"4d",x"10",x"30",x"4d",x"10",x"1f",x"02",x"8d",x"10",x"1f",x"11",x"15",x"12",x"34",x"cd",x"10",x"1f",x"11",x"15",x"15",x"00",x"f2",x"7b",x"00",x"25",x"60",x"10",x"10",x"5f",x"15",x"42",x"10",x"7b",x"00",x"e9",x"55",x"00",x"c0",x"c1",x"6d",x"10",x"40",x"f5",x"e0",x"10",x"5e",x"15",x"22",x"10",x"5e",x"15",x"12",x"10",x"00",x"20",x"10",x"5e",x"15",x"02",x"63",x"11",x"60",x"10",x"00",x"64",x"00",x"5c",x"01",x"00",x"60",x"5d",x"03",x"08",x"2f",x"a2",x"12",x"00",x"54",x"5e",x"02",x"00",x"58",x"00",x"48",x"00",x"44",x"08",x"2f",x"61",x"12",x"01",x"40",x"25",x"21",x"80",x"10",x"40",x"35",x"08",x"1f",x"41",x"43",x"00",x"51",x"62",x"14",x"15",x"11",x"40",x"20",x"23",x"20",x"10",x"3c",x"00",x"54",x"43",x"00",x"41",x"62",x"14",x"15",x"11",x"40",x"20",x"32",x"e0",x"10",x"3e",x"00",x"58",x"43",x"00",x"51",x"62",x"14",x"15",x"11",x"40",x"00",x"44",x"00",x"48",x"12",x"00",x"12",x"01",x"11",x"20",x"10",x"00",x"5c",x"00",x"60",x"00",x"64",x"00",x"44",x"00",x"64",x"00",x"60",x"00",x"5c",x"13",x"08",x"1f",x"51",x"2f",x"ed",x"10",x"5f",x"2d",x"10",x"0d",x"10",x"51",x"c3",x"13",x"41",x"2d",x"c2",x"04",x"08",x"2f",x"4d",x"10",x"01",x"00",x"05",x"00",x"50",x"03",x"4d",x"10",x"11",x"00",x"01",x"08",x"5f",x"12",x"01",x"00",x"01",x"2f",x"11",x"01",x"44",x"14",x"c6",x"2d",x"13",x"62",x"8d",x"10",x"c1",x"c3",x"12",x"51",x"2c",x"c2",x"80",x"04",x"08",x"2f",x"4d",x"10",x"01",x"00",x"05",x"00",x"50",x"00",x"03",x"0d",x"10",x"11",x"00",x"01",x"00",x"44",x"00",x"48",x"00",x"64",x"23",x"12",x"01",x"00",x"31",x"ad",x"10",x"05",x"2f",x"15",x"02",x"60",x"12",x"91",x"02",x"2d",x"10",x"60",x"60",x"12",x"d1",x"42",x"6d",x"10",x"61",x"ad",x"10",x"50",x"12",x"e0",x"10",x"00",x"44",x"10",x"00",x"44",x"02",x"00",x"08",x"4f",x"02",x"63",x"41",x"01",x"31",x"51",x"6d",x"10",x"ff",x"f1",x"02",x"12",x"ff",x"1f",x"05",x"22",x"02",x"00",x"25",x"20",x"10",x"00",x"4c",x"06",x"05",x"21",x"41",x"3c",x"61",x"11",x"15",x"00",x"15",x"16",x"60",x"10",x"50",x"12",x"63",x"11",x"00",x"4c",x"00",x"01",x"00",x"02",x"63",x"41",x"21",x"71",x"3e",x"61",x"10",x"15",x"00",x"67",x"02",x"12",x"ff",x"01",x"00",x"02",x"63",x"41",x"21",x"71",x"38",x"61",x"10",x"15",x"00",x"47",x"02",x"12",x"ff",x"08",x"2f",x"ff",x"f1",x"01",x"00",x"60",x"21",x"a0",x"10",x"61",x"00",x"51",x"ed",x"10",x"00",x"60",x"00",x"10",x"63",x"4c",x"21",x"4d",x"10",x"08",x"1f",x"c5",x"2a",x"13",x"52",x"4d",x"10",x"01",x"c3",x"60",x"04",x"61",x"0f",x"91",x"42",x"2d",x"10",x"60",x"10",x"62",x"0f",x"08",x"1f",x"cd",x"10",x"1c",x"20",x"24",x"01",x"08",x"10",x"0f",x"4f",x"5f",x"35",x"0c",x"08",x"04",x"2f",x"72",x"10",x"cd",x"10",x"08",x"0c",x"0f",x"10",x"9f",x"df",x"0c",x"08",x"2e",x"04",x"60",x"10",x"f0",x"1f",x"01",x"02",x"2a",x"1a",x"77",x"37",x"98",x"80",x"10",x"51",x"ff",x"01",x"02",x"2a",x"1a",x"87",x"88",x"38",x"88",x"89",x"87",x"ff",x"11",x"e0",x"10",x"14",x"02",x"03",x"07",x"78",x"99",x"e9",x"bf",x"93",x"a0",x"10",x"03",x"10",x"a9",x"00",x"0b",x"18",x"58",x"ff",x"11",x"51",x"ff",x"21",x"e6",x"0e",x"bf",x"6e",x"12",x"02",x"07",x"08",x"01",x"0a",x"01",x"58",x"01",x"ba",x"aa",x"aa",x"09",x"a0",x"10",x"31",x"e0",x"10",x"03",x"07",x"08",x"89",x"aa",x"ea",x"6f",x"a7",x"a0",x"10",x"07",x"10",x"1e",x"40",x"10",x"e3",x"19",x"59",x"ff",x"11",x"51",x"ff",x"31",x"8d",x"10",x"05",x"01",x"2f",x"01",x"2f",x"15",x"07",x"08",x"09",x"88",x"e8",x"a5",x"3a",x"1a",x"7e",x"01",x"01",x"4e",x"ee",x"ee",x"0b",x"40",x"10",x"6e",x"57",x"ff",x"11",x"40",x"10",x"10",x"03",x"07",x"08",x"89",x"aa",x"ea",x"a7",x"a0",x"10",x"07",x"10",x"1e",x"40",x"10",x"e3",x"19",x"59",x"ff",x"11",x"51",x"ff",x"2f",x"31",x"cd",x"10",x"05",x"01",x"6e",x"20",x"f3",x"ef",x"6f",x"15",x"09",x"1c",x"01",x"11",x"1e",x"0e",x"8e",x"11",x"61",x"12",x"01",x"5e",x"11",x"41",x"11",x"02",x"05",x"02",x"72",x"01",x"40",x"10",x"19",x"18",x"20",x"10",x"1c",x"51",x"ff",x"01",x"0a",x"15",x"08",x"02",x"02",x"92",x"10",x"23",x"00",x"a4",x"00",x"1b",x"40",x"10",x"b4",x"9a",x"60",x"10",x"9a",x"40",x"10",x"20",x"10",x"02",x"14",x"0b",x"12",x"0d",x"10",x"01",x"4d",x"10",x"41",x"0b",x"05",x"00",x"af",x"bf",x"02",x"03",x"37",x"17",x"88",x"b8",x"a9",x"98",x"ff",x"12",x"60",x"10",x"10",x"0d",x"10",x"04",x"08",x"0c",x"11",x"d0",x"01",x"00",x"07",x"08",x"89",x"19",x"aa",x"2a",x"3b",x"80",x"10",x"17",x"ff",x"d0",x"00",x"4f",x"80",x"10",x"71",x"09",x"0b",x"19",x"02",x"01",x"2a",x"bb",x"0b",x"e0",x"10",x"17",x"ff",x"4f",x"d0",x"8f",x"4f",x"5f",x"40",x"10",x"07",x"09",x"0a",x"ab",x"ee",x"2e",x"e9",x"a0",x"10",x"09",x"10",x"4e",x"00",x"05",x"1b",x"1b",x"ff",x"18",x"18",x"ff",x"5f",x"04",x"8f",x"10",x"4f",x"5f",x"80",x"10",x"78",x"71",x"09",x"28",x"ab",x"be",x"1b",x"55",x"4e",x"ee",x"ee",x"e5",x"e9",x"ff",x"17",x"17",x"ff",x"5f",x"04",x"d0",x"4f",x"08",x"04",x"01",x"00",x"07",x"08",x"89",x"0b",x"aa",x"2a",x"e1",x"8e",x"1e",x"96",x"01",x"01",x"46",x"66",x"66",x"05",x"40",x"10",x"ba",x"80",x"10",x"17",x"ff",x"6f",x"04",x"08",x"d0",x"cf",x"08",x"04",x"2f",x"01",x"00",x"07",x"f9",x"0a",x"7f",x"8f",x"ab",x"05",x"77",x"78",x"0e",x"08",x"07",x"16",x"77",x"88",x"37",x"77",x"77",x"87",x"78",x"77",x"28",x"78",x"75",x"ff",x"1b",x"1b",x"ff",x"7f",x"17",x"a0",x"10",x"5f",x"4f",x"4f",x"10",x"0f",x"18",x"08",x"04",x"4f",x"03",x"00",x"38",x"07",x"00",x"03",x"13",x"33",x"99",x"79",x"ff",x"32",x"01",x"11",x"60",x"10",x"09",x"0e",x"76",x"08",x"ff",x"8a",x"aa",x"8a",x"a8",x"e5",x"15",x"3a",x"aa",x"bb",x"2a",x"04",x"0b",x"6b",x"00",x"b4",x"60",x"10",x"17",x"20",x"10",x"0c",x"01",x"02",x"28",x"32",x"08",x"0c",x"6f",x"04",x"08",x"d0",x"4f",x"4f",x"5f",x"25",x"04",x"54",x"4c",x"48",x"44",x"40",x"3c",x"38",x"34",x"2c",x"28",x"24",x"20",x"1c",x"18",x"14",x"30",x"10",x"36",x"50",x"01",x"00",x"20",x"f1",x"f2",x"8d",x"10",x"02",x"10",x"21",x"21",x"50",x"01",x"00",x"20",x"3f",x"41",x"50",x"15",x"1f",x"00",x"10",x"21",x"60",x"10",x"21",x"41",x"ff",x"1f",x"5f",x"36",x"01",x"00",x"20",x"f1",x"f2",x"cd",x"10",x"02",x"10",x"21",x"21",x"50",x"01",x"00",x"20",x"5f",x"1f",x"11",x"00",x"2f",x"15",x"60",x"10",x"15",x"45",x"ff",x"5f",x"2f",x"1f",x"6d",x"10",x"1f",x"ad",x"10",x"1f",x"ed",x"10",x"1f",x"2d",x"10",x"1f",x"6d",x"10",x"1f",x"ad",x"10",x"1f",x"ed",x"10",x"1f",x"2d",x"10",x"1f",x"6d",x"10",x"1f",x"ad",x"10",x"1f",x"ed",x"10",x"1f",x"2d",x"10",x"1f",x"6d",x"10",x"1f",x"ad",x"10",x"1f",x"ed",x"10",x"1f",x"2d",x"10",x"04",x"08",x"0c",x"cf",x"10",x"71",x"a7",x"80",x"10",x"01",x"03",x"00",x"8a",x"cb",x"00",x"00",x"10",x"80",x"10",x"00",x"10",x"80",x"10",x"00",x"a3",x"83",x"80",x"10",x"08",x"32",x"43",x"01",x"53",x"00",x"43",x"00",x"a0",x"10",x"20",x"10",x"10",x"32",x"53",x"01",x"63",x"00",x"80",x"10",x"18",x"32",x"a3",x"83",x"73",x"40",x"10",x"00",x"a3",x"83",x"43",x"60",x"10",x"bb",x"00",x"db",x"00",x"eb",x"00",x"53",x"00",x"33",x"00",x"bb",x"00",x"db",x"00",x"32",x"13",x"0c",x"00",x"10",x"80",x"10",x"03",x"53",x"00",x"32",x"13",x"14",x"a0",x"73",x"00",x"a3",x"83",x"73",x"00",x"10",x"00",x"32",x"eb",x"32",x"53",x"00",x"13",x"10",x"d0",x"0a",x"aa",x"00",x"60",x"a3",x"83",x"53",x"80",x"10",x"10",x"04",x"32",x"13",x"1a",x"a7",x"7b",x"0a",x"00",x"b7",x"c0",x"10",x"10",x"60",x"7b",x"b1",x"d0",x"32",x"13",x"0c",x"10",x"04",x"32",x"a0",x"32",x"13",x"10",x"10",x"14",x"32",x"7b",x"13",x"10",x"df",x"0c",x"08",x"04",x"10",x"ff",x"c9",x"0e",x"10",x"0b",x"eb",x"a1",x"17",x"5b",x"8b",x"00",x"a0",x"10",x"01",x"00",x"76",x"6e",x"16",x"3b",x"ab",x"ff",x"47",x"0a",x"12",x"25",x"06",x"a0",x"10",x"a0",x"10",x"fd",x"c0",x"10",x"10",x"fb",x"c0",x"10",x"40",x"10",x"01",x"a1",x"5e",x"ff",x"51",x"ca",x"0a",x"20",x"10",x"01",x"a1",x"5e",x"0b",x"eb",x"ff",x"51",x"ca",x"0a",x"60",x"10",x"10",x"40",x"10",x"02",x"03",x"02",x"1d",x"6f",x"5f",x"4f",x"df",x"d0",x"12",x"22",x"00",x"12",x"00",x"60",x"41",x"20",x"32",x"00",x"42",x"00",x"20",x"c1",x"60",x"22",x"00",x"81",x"60",x"81",x"e0",x"52",x"00",x"c1",x"11",x"10",x"40",x"08",x"78",x"09",x"00",x"32",x"01",x"0f",x"89",x"01",x"02",x"40",x"10",x"ff",x"e2",x"0f",x"9a",x"8a",x"18",x"a8",x"0a",x"40",x"10",x"29",x"0f",x"01",x"09",x"03",x"78",x"0a",x"00",x"39",x"88",x"9a",x"8a",x"18",x"a8",x"0a",x"40",x"10",x"29",x"0f",x"01",x"09",x"05",x"78",x"0a",x"00",x"39",x"88",x"9a",x"8a",x"18",x"a8",x"0a",x"40",x"10",x"29",x"07",x"01",x"71",x"87",x"0a",x"40",x"10",x"72",x"0f",x"01",x"ff",x"f2",x"d0",x"8f",x"4f",x"14",x"00",x"ed",x"10",x"41",x"2d",x"10",x"04",x"8f",x"10",x"df",x"08",x"04",x"f5",x"54",x"ad",x"10",x"ff",x"01",x"11",x"6d",x"10",x"41",x"51",x"fe",x"12",x"18",x"fe",x"5f",x"4f",x"df",x"d0",x"8f",x"4f",x"14",x"00",x"6d",x"10",x"ff",x"01",x"11",x"2d",x"10",x"04",x"8f",x"10",x"d0",x"23",x"04",x"07",x"ff",x"21",x"10",x"63",x"22",x"04",x"07",x"ff",x"12",x"10",x"fd",x"4f",x"5f",x"6f",x"02",x"4f",x"02",x"3f",x"02",x"2f",x"24",x"f2",x"00",x"01",x"2f",x"00",x"2f",x"88",x"f2",x"00",x"00",x"02",x"2f",x"60",x"61",x"21",x"c0",x"10",x"87",x"00",x"18",x"10",x"21",x"01",x"01",x"a3",x"00",x"03",x"00",x"60",x"7b",x"c0",x"b3",x"00",x"03",x"00",x"e0",x"8b",x"00",x"33",x"00",x"01",x"10",x"80",x"d3",x"00",x"01",x"10",x"d0",x"97",x"80",x"10",x"01",x"08",x"12",x"38",x"17",x"13",x"a7",x"ff",x"00",x"f8",x"a3",x"00",x"00",x"2f",x"c3",x"32",x"04",x"00",x"d8",x"12",x"f8",x"00",x"01",x"01",x"08",x"f1",x"60",x"10",x"10",x"00",x"f4",x"00",x"e8",x"01",x"01",x"d0",x"08",x"98",x"00",x"32",x"01",x"07",x"1b",x"27",x"38",x"32",x"a8",x"ff",x"20",x"01",x"bf",x"01",x"8f",x"01",x"2f",x"f6",x"10",x"93",x"a8",x"00",x"00",x"3f",x"c7",x"02",x"73",x"04",x"00",x"d8",x"32",x"06",x"00",x"e4",x"40",x"10",x"02",x"92",x"60",x"10",x"10",x"00",x"e4",x"01",x"01",x"1f",x"31",x"10",x"27",x"87",x"00",x"27",x"00",x"17",x"00",x"87",x"00",x"00",x"10",x"00",x"f4",x"12",x"00",x"f4",x"10",x"c0",x"10",x"c0",x"10",x"80",x"10",x"03",x"83",x"10",x"a0",x"10",x"80",x"10",x"04",x"01",x"2f",x"21",x"01",x"2f",x"20",x"37",x"04",x"57",x"00",x"87",x"00",x"80",x"10",x"00",x"1f",x"c2",x"21",x"04",x"00",x"d8",x"01",x"1f",x"1f",x"6f",x"51",x"00",x"e8",x"0f",x"15",x"00",x"e4",x"fd",x"01",x"3f",x"02",x"01",x"3f",x"00",x"17",x"00",x"40",x"10",x"00",x"f0",x"06",x"00",x"2f",x"32",x"23",x"00",x"3f",x"03",x"01",x"2f",x"80",x"10",x"01",x"01",x"af",x"01",x"6f",x"01",x"62",x"01",x"00",x"f2",x"01",x"bf",x"f8",x"1b",x"03",x"04",x"21",x"11",x"18",x"19",x"1a",x"01",x"04",x"27",x"77",x"1b",x"3f",x"9f",x"3b",x"37",x"83",x"23",x"7f",x"33",x"1f",x"20",x"03",x"04",x"27",x"77",x"21",x"3f",x"9f",x"3b",x"37",x"83",x"23",x"7f",x"33",x"25",x"26",x"05",x"04",x"27",x"77",x"27",x"2f",x"02",x"00",x"f0",x"02",x"00",x"40",x"10",x"00",x"e8",x"80",x"10",x"06",x"f4",x"02",x"0d",x"10",x"18",x"04",x"05",x"03",x"00",x"67",x"10",x"18",x"67",x"61",x"01",x"1f",x"01",x"3f",x"31",x"04",x"00",x"f1",x"02",x"20",x"10",x"c0",x"10",x"18",x"01",x"7f",x"71",x"41",x"33",x"a6",x"42",x"11",x"41",x"34",x"a2",x"8d",x"10",x"a2",x"15",x"41",x"34",x"01",x"7f",x"14",x"00",x"a4",x"00",x"00",x"f1",x"a2",x"00",x"e0",x"05",x"0d",x"10",x"62",x"61",x"15",x"cd",x"10",x"00",x"e0",x"17",x"10",x"62",x"00",x"18",x"71",x"22",x"01",x"3f",x"76",x"13",x"40",x"10",x"00",x"f4",x"21",x"80",x"10",x"02",x"01",x"2f",x"01",x"5f",x"21",x"26",x"00",x"60",x"10",x"04",x"02",x"00",x"e0",x"0d",x"10",x"00",x"e0",x"01",x"7f",x"e0",x"10",x"80",x"10",x"00",x"d8",x"31",x"12",x"00",x"2f",x"01",x"3f",x"12",x"40",x"10",x"01",x"3f",x"84",x"21",x"08",x"04",x"00",x"01",x"4f",x"51",x"2d",x"10",x"a0",x"10",x"00",x"f4",x"21",x"80",x"10",x"01",x"01",x"6f",x"01",x"1f",x"64",x"14",x"00",x"c0",x"10",x"02",x"4d",x"10",x"00",x"d8",x"31",x"12",x"00",x"2f",x"45",x"65",x"12",x"04",x"67",x"00",x"00",x"1f",x"82",x"71",x"42",x"00",x"2f",x"11",x"00",x"e0",x"00",x"d8",x"04",x"00",x"d8",x"00",x"f4",x"73",x"02",x"00",x"40",x"10",x"01",x"5f",x"23",x"01",x"51",x"52",x"00",x"01",x"2f",x"a0",x"10",x"00",x"d8",x"31",x"12",x"00",x"2f",x"81",x"60",x"10",x"62",x"84",x"a0",x"10",x"84",x"e0",x"10",x"01",x"01",x"e0",x"10",x"41",x"60",x"10",x"00",x"f4",x"84",x"21",x"c0",x"10",x"00",x"e8",x"80",x"10",x"02",x"81",x"41",x"51",x"00",x"ec",x"00",x"e0",x"11",x"01",x"8f",x"f1",x"41",x"00",x"e8",x"00",x"ec",x"00",x"10",x"15",x"01",x"2f",x"12",x"60",x"10",x"10",x"ff",x"c0",x"10",x"15",x"01",x"f7",x"02",x"09",x"25",x"11",x"f7",x"01",x"6f",x"01",x"4f",x"00",x"01",x"4f",x"80",x"10",x"00",x"f0",x"02",x"16",x"00",x"d8",x"43",x"13",x"21",x"04",x"00",x"d8",x"15",x"01",x"02",x"15",x"01",x"f7",x"01",x"5f",x"32",x"01",x"3f",x"03",x"01",x"2f",x"21",x"00",x"ec",x"00",x"e0",x"1b",x"15",x"40",x"10",x"01",x"2f",x"01",x"04",x"01",x"1f",x"01",x"1f",x"01",x"2f",x"cd",x"10",x"11",x"00",x"01",x"00",x"f8",x"51",x"02",x"2f",x"12",x"01",x"2f",x"01",x"01",x"8f",x"82",x"00",x"01",x"2f",x"00",x"01",x"f7",x"12",x"00",x"e0",x"00",x"e8",x"20",x"10",x"f7",x"81",x"80",x"10",x"01",x"81",x"03",x"1f",x"28",x"01",x"2f",x"11",x"12",x"60",x"10",x"01",x"1f",x"16",x"00",x"18",x"83",x"15",x"80",x"10",x"01",x"13",x"01",x"61",x"ff",x"65",x"00",x"e8",x"16",x"f8",x"48",x"21",x"00",x"10",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"1f",x"15",x"51",x"60",x"10",x"10",x"ef",x"a0",x"10",x"61",x"80",x"10",x"00",x"e8",x"52",x"60",x"10",x"18",x"11",x"33",x"12",x"ff",x"61",x"40",x"10",x"15",x"00",x"e8",x"16",x"f7",x"f1",x"12",x"51",x"43",x"0e",x"45",x"00",x"e4",x"80",x"10",x"00",x"e8",x"f1",x"06",x"00",x"62",x"00",x"0c",x"08",x"71",x"91",x"00",x"91",x"18",x"25",x"00",x"14",x"00",x"10",x"00",x"e8",x"60",x"10",x"f5",x"61",x"00",x"f8",x"04",x"02",x"4f",x"71",x"01",x"f1",x"f4",x"1f",x"f1",x"1f",x"01",x"1f",x"01",x"2f",x"01",x"6f",x"63",x"0c",x"1f",x"62",x"a0",x"10",x"40",x"10",x"ff",x"38",x"00",x"f8",x"01",x"30",x"08",x"34",x"04",x"00",x"fc",x"00",x"e0",x"00",x"ec",x"0c",x"2f",x"02",x"00",x"88",x"f2",x"10",x"00",x"2f",x"02",x"2f",x"31",x"32",x"00",x"14",x"00",x"00",x"e3",x"02",x"01",x"10",x"01",x"00",x"10",x"00",x"fc",x"12",x"71",x"73",x"21",x"ff",x"51",x"40",x"10",x"56",x"02",x"2f",x"12",x"30",x"c0",x"10",x"00",x"e0",x"00",x"ec",x"04",x"19",x"f4",x"c0",x"10",x"60",x"14",x"03",x"02",x"01",x"1f",x"80",x"10",x"00",x"fc",x"43",x"61",x"00",x"01",x"1f",x"b2",x"21",x"a2",x"24",x"02",x"5f",x"01",x"15",x"41",x"22",x"a2",x"23",x"01",x"15",x"01",x"1f",x"16",x"4d",x"10",x"cd",x"10",x"54",x"f5",x"16",x"01",x"01",x"2f",x"02",x"9f",x"21",x"00",x"f8",x"40",x"10",x"02",x"2f",x"40",x"10",x"10",x"72",x"60",x"10",x"40",x"10",x"40",x"10",x"10",x"01",x"a0",x"10",x"e0",x"10",x"78",x"77",x"07",x"00",x"f3",x"03",x"ff",x"28",x"13",x"00",x"32",x"f3",x"87",x"01",x"ff",x"60",x"82",x"e3",x"59",x"72",x"00",x"01",x"00",x"01",x"00",x"18",x"13",x"40",x"10",x"11",x"e7",x"00",x"83",x"e0",x"10",x"07",x"00",x"60",x"13",x"72",x"20",x"10",x"a0",x"10",x"40",x"10",x"78",x"ff",x"ff",x"00",x"10",x"60",x"10",x"fe",x"e0",x"10",x"88",x"f2",x"01",x"03",x"01",x"cd",x"10",x"00",x"88",x"00",x"f4",x"00",x"0c",x"00",x"03",x"27",x"21",x"00",x"71",x"77",x"07",x"00",x"f3",x"03",x"ff",x"21",x"12",x"04",x"02",x"00",x"14",x"00",x"a0",x"88",x"f2",x"00",x"f0",x"12",x"02",x"43",x"0a",x"01",x"8f",x"46",x"01",x"6f",x"40",x"f4",x"00",x"e8",x"00",x"01",x"00",x"01",x"1f",x"21",x"01",x"1f",x"01",x"01",x"00",x"14",x"00",x"20",x"02",x"2f",x"01",x"6f",x"f1",x"43",x"61",x"09",x"46",x"01",x"6f",x"40",x"f4",x"00",x"e4",x"00",x"f0",x"05",x"00",x"01",x"5f",x"a0",x"12",x"00",x"13",x"51",x"32",x"00",x"60",x"01",x"1f",x"51",x"14",x"ef",x"51",x"43",x"09",x"45",x"01",x"ef",x"12",x"f1",x"f4",x"63",x"08",x"34",x"04",x"00",x"e0",x"00",x"ec",x"08",x"2f",x"02",x"00",x"88",x"f4",x"10",x"00",x"2f",x"02",x"4f",x"31",x"60",x"10",x"10",x"16",x"80",x"10",x"00",x"e1",x"63",x"01",x"02",x"08",x"46",x"14",x"60",x"10",x"30",x"07",x"00",x"e2",x"07",x"24",x"84",x"02",x"00",x"80",x"84",x"12",x"30",x"03",x"c0",x"10",x"02",x"fc",x"24",x"01",x"21",x"31",x"60",x"10",x"10",x"30",x"11",x"a0",x"10",x"34",x"31",x"14",x"01",x"a0",x"10",x"10",x"e0",x"10",x"15",x"00",x"dc",x"60",x"10",x"00",x"43",x"27",x"a9",x"7a",x"40",x"10",x"11",x"89",x"28",x"98",x"a0",x"10",x"0c",x"10",x"14",x"cf",x"d0",x"00",x"df",x"0c",x"08",x"04",x"29",x"1f",x"17",x"02",x"00",x"e2",x"07",x"aa",x"21",x"60",x"10",x"63",x"32",x"22",x"02",x"21",x"71",x"80",x"10",x"60",x"10",x"10",x"71",x"80",x"10",x"b2",x"10",x"f4",x"91",x"a0",x"71",x"02",x"1f",x"81",x"11",x"14",x"01",x"64",x"08",x"8f",x"60",x"10",x"10",x"60",x"10",x"10",x"2f",x"80",x"2f",x"00",x"2f",x"03",x"00",x"e4",x"72",x"03",x"68",x"60",x"32",x"1f",x"80",x"10",x"54",x"58",x"10",x"95",x"1f",x"91",x"26",x"2f",x"21",x"2f",x"12",x"42",x"24",x"19",x"09",x"ff",x"c0",x"01",x"54",x"10",x"58",x"1f",x"16",x"00",x"16",x"54",x"68",x"60",x"64",x"03",x"21",x"40",x"10",x"60",x"10",x"10",x"02",x"0d",x"10",x"f3",x"10",x"2f",x"f1",x"21",x"60",x"10",x"14",x"70",x"01",x"00",x"05",x"00",x"20",x"81",x"01",x"14",x"00",x"85",x"00",x"01",x"14",x"60",x"58",x"21",x"e0",x"10",x"60",x"10",x"10",x"6c",x"00",x"76",x"41",x"05",x"64",x"40",x"f7",x"54",x"00",x"10",x"51",x"02",x"61",x"8d",x"10",x"5f",x"46",x"05",x"00",x"51",x"f1",x"10",x"13",x"32",x"c0",x"10",x"17",x"00",x"80",x"41",x"73",x"0d",x"10",x"01",x"10",x"6f",x"5f",x"4f",x"df",x"d0",x"cf",x"df",x"10",x"0c",x"63",x"08",x"18",x"04",x"10",x"10",x"4f",x"10",x"df",x"0c",x"08",x"04",x"28",x"03",x"2f",x"1f",x"0d",x"10",x"01",x"00",x"06",x"24",x"20",x"04",x"0e",x"f1",x"40",x"10",x"2f",x"61",x"02",x"00",x"27",x"e7",x"03",x"24",x"40",x"10",x"2f",x"2f",x"03",x"e0",x"10",x"32",x"00",x"21",x"20",x"10",x"04",x"1f",x"cf",x"03",x"06",x"10",x"24",x"14",x"2c",x"0f",x"01",x"00",x"1f",x"03",x"50",x"38",x"24",x"2c",x"20",x"80",x"04",x"12",x"f3",x"c2",x"04",x"c2",x"7f",x"1e",x"84",x"1c",x"18",x"04",x"c2",x"80",x"04",x"1b",x"c2",x"19",x"01",x"04",x"ff",x"10",x"24",x"14",x"2c",x"10",x"2f",x"3f",x"01",x"24",x"13",x"ff",x"7f",x"76",x"00",x"40",x"10",x"44",x"26",x"28",x"76",x"ff",x"7f",x"2f",x"c0",x"10",x"28",x"30",x"04",x"0d",x"01",x"40",x"10",x"1f",x"03",x"1f",x"2f",x"cd",x"10",x"11",x"00",x"01",x"20",x"12",x"01",x"00",x"60",x"2f",x"1f",x"00",x"03",x"6f",x"2f",x"1f",x"cd",x"10",x"00",x"03",x"1f",x"62",x"0e",x"3f",x"01",x"28",x"36",x"c0",x"10",x"18",x"44",x"1c",x"24",x"2c",x"e0",x"7f",x"2f",x"c0",x"7f",x"2f",x"03",x"44",x"24",x"48",x"24",x"02",x"00",x"03",x"34",x"02",x"00",x"21",x"2f",x"78",x"20",x"00",x"1f",x"01",x"1f",x"80",x"10",x"24",x"00",x"03",x"86",x"19",x"f3",x"c2",x"02",x"1f",x"c4",x"18",x"1c",x"17",x"7f",x"01",x"18",x"78",x"00",x"1f",x"18",x"ff",x"1f",x"01",x"00",x"40",x"17",x"48",x"12",x"7a",x"17",x"44",x"10",x"21",x"10",x"44",x"21",x"c0",x"73",x"17",x"ff",x"73",x"a7",x"00",x"83",x"60",x"10",x"10",x"09",x"17",x"80",x"10",x"40",x"10",x"1a",x"10",x"2a",x"04",x"08",x"0c",x"cf",x"10",x"cf",x"df",x"10",x"0c",x"1c",x"08",x"18",x"04",x"fc",x"4f",x"df",x"d0",x"00",x"47",x"df",x"10",x"0c",x"08",x"18",x"04",x"fb",x"4f",x"df",x"d0",x"00",x"7f",x"df",x"10",x"0c",x"08",x"18",x"04",x"fb",x"4f",x"df",x"d0",x"d0",x"d0",x"d0",x"01",x"10",x"8f",x"4f",x"8d",x"10",x"e3",x"03",x"8d",x"10",x"04",x"8f",x"10",x"12",x"d0",x"02",x"d0",x"38",x"07",x"60",x"10",x"10",x"03",x"00",x"27",x"f3",x"09",x"80",x"10",x"10",x"43",x"00",x"f8",x"f3",x"89",x"98",x"10",x"00",x"10",x"87",x"87",x"87",x"03",x"f3",x"ff",x"80",x"87",x"c3",x"40",x"10",x"00",x"10",x"f3",x"03",x"ff",x"d0",x"8f",x"14",x"07",x"4f",x"87",x"ff",x"38",x"00",x"f8",x"00",x"00",x"10",x"00",x"87",x"17",x"28",x"60",x"10",x"10",x"04",x"17",x"03",x"73",x"10",x"40",x"10",x"ff",x"f7",x"08",x"09",x"c0",x"10",x"13",x"04",x"04",x"cd",x"10",x"40",x"13",x"04",x"00",x"21",x"00",x"00",x"07",x"73",x"04",x"04",x"2c",x"d0",x"4f",x"4f",x"5f",x"25",x"1a",x"ff",x"6f",x"75",x"1a",x"72",x"17",x"ff",x"18",x"00",x"08",x"19",x"00",x"09",x"00",x"89",x"08",x"07",x"c0",x"10",x"14",x"17",x"11",x"ff",x"18",x"00",x"08",x"19",x"00",x"09",x"00",x"89",x"01",x"01",x"11",x"05",x"00",x"08",x"00",x"02",x"00",x"09",x"00",x"98",x"01",x"00",x"00",x"01",x"a1",x"00",x"10",x"18",x"40",x"10",x"19",x"ff",x"40",x"10",x"40",x"10",x"81",x"40",x"10",x"00",x"48",x"8c",x"05",x"00",x"01",x"08",x"08",x"00",x"3a",x"00",x"03",x"01",x"12",x"ff",x"02",x"00",x"a1",x"40",x"10",x"2c",x"05",x"71",x"01",x"00",x"48",x"8c",x"05",x"25",x"01",x"00",x"60",x"10",x"01",x"01",x"a0",x"10",x"18",x"40",x"10",x"27",x"00",x"01",x"00",x"18",x"08",x"00",x"57",x"00",x"45",x"40",x"10",x"40",x"10",x"f3",x"21",x"a6",x"09",x"00",x"09",x"08",x"00",x"2f",x"00",x"10",x"1c",x"60",x"10",x"01",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"18",x"10",x"01",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"11",x"21",x"43",x"81",x"cd",x"10",x"c1",x"41",x"61",x"f2",x"6f",x"21",x"ff",x"f1",x"61",x"00",x"8f",x"7f",x"a0",x"10",x"18",x"c0",x"10",x"01",x"14",x"12",x"02",x"23",x"32",x"08",x"23",x"32",x"32",x"aa",x"27",x"73",x"02",x"66",x"32",x"22",x"32",x"23",x"32",x"1e",x"32",x"02",x"23",x"24",x"e0",x"52",x"96",x"14",x"23",x"32",x"04",x"23",x"32",x"10",x"f3",x"55",x"53",x"01",x"32",x"33",x"33",x"07",x"02",x"72",x"04",x"0f",x"f3",x"01",x"13",x"02",x"22",x"32",x"43",x"52",x"03",x"c2",x"69",x"0a",x"03",x"1d",x"03",x"31",x"01",x"31",x"a0",x"10",x"21",x"10",x"05",x"06",x"60",x"10",x"53",x"10",x"28",x"11",x"cf",x"16",x"2f",x"51",x"41",x"02",x"1c",x"11",x"40",x"10",x"2f",x"9f",x"21",x"20",x"1c",x"07",x"00",x"f7",x"2f",x"2f",x"8f",x"22",x"83",x"23",x"03",x"01",x"83",x"00",x"a0",x"21",x"36",x"00",x"03",x"03",x"01",x"47",x"53",x"21",x"44",x"19",x"21",x"05",x"01",x"25",x"63",x"15",x"31",x"01",x"02",x"01",x"ff",x"f4",x"01",x"9f",x"04",x"00",x"41",x"41",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"11",x"60",x"10",x"01",x"01",x"60",x"10",x"08",x"01",x"80",x"10",x"01",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"11",x"21",x"f8",x"52",x"8d",x"10",x"10",x"c5",x"09",x"07",x"00",x"2f",x"00",x"01",x"8c",x"80",x"10",x"e0",x"10",x"01",x"02",x"03",x"2f",x"52",x"00",x"c1",x"40",x"10",x"3f",x"41",x"8d",x"10",x"c6",x"09",x"03",x"00",x"53",x"07",x"12",x"1d",x"03",x"3f",x"32",x"14",x"73",x"43",x"00",x"08",x"72",x"43",x"00",x"12",x"82",x"31",x"6f",x"5f",x"4f",x"df",x"d0",x"07",x"07",x"00",x"31",x"03",x"01",x"00",x"03",x"00",x"07",x"01",x"07",x"07",x"02",x"71",x"2c",x"10",x"cf",x"1a",x"02",x"00",x"0a",x"ff",x"1b",x"08",x"ff",x"40",x"10",x"40",x"10",x"7a",x"80",x"10",x"1a",x"04",x"00",x"0b",x"00",x"09",x"00",x"0e",x"00",x"eb",x"0a",x"00",x"89",x"24",x"78",x"08",x"00",x"13",x"07",x"00",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"20",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"98",x"f7",x"40",x"10",x"31",x"21",x"40",x"10",x"4f",x"4f",x"10",x"cf",x"1a",x"02",x"00",x"0a",x"ff",x"1b",x"08",x"ff",x"40",x"10",x"40",x"10",x"7a",x"0a",x"00",x"39",x"1b",x"40",x"10",x"1e",x"ff",x"40",x"10",x"40",x"10",x"ba",x"60",x"10",x"07",x"08",x"07",x"20",x"10",x"07",x"60",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"80",x"10",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"40",x"10",x"87",x"f7",x"00",x"17",x"42",x"01",x"00",x"07",x"71",x"d0",x"cf",x"ff",x"02",x"4f",x"11",x"00",x"02",x"ff",x"17",x"00",x"07",x"00",x"72",x"02",x"00",x"ff",x"f1",x"04",x"11",x"00",x"01",x"ff",x"40",x"10",x"40",x"10",x"4f",x"d0",x"00",x"17",x"4f",x"40",x"10",x"ff",x"f9",x"91",x"00",x"08",x"00",x"0b",x"00",x"ba",x"0a",x"00",x"39",x"1b",x"40",x"10",x"1e",x"ff",x"40",x"10",x"40",x"10",x"ba",x"60",x"10",x"07",x"08",x"07",x"20",x"10",x"07",x"60",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"80",x"10",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"40",x"10",x"78",x"08",x"00",x"17",x"42",x"01",x"00",x"07",x"71",x"d0",x"00",x"17",x"4f",x"40",x"10",x"ff",x"f9",x"91",x"00",x"08",x"00",x"0b",x"00",x"ba",x"0a",x"00",x"39",x"1b",x"40",x"10",x"1e",x"ff",x"40",x"10",x"40",x"10",x"ba",x"60",x"10",x"07",x"08",x"07",x"20",x"10",x"07",x"60",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"80",x"10",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"40",x"10",x"78",x"08",x"00",x"17",x"42",x"01",x"00",x"07",x"71",x"d0",x"00",x"17",x"4f",x"40",x"10",x"ff",x"f9",x"91",x"00",x"08",x"00",x"0b",x"00",x"ba",x"0a",x"00",x"39",x"1b",x"40",x"10",x"1e",x"ff",x"40",x"10",x"40",x"10",x"ba",x"60",x"10",x"07",x"08",x"07",x"20",x"10",x"07",x"60",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"80",x"10",x"10",x"18",x"40",x"10",x"19",x"40",x"10",x"40",x"10",x"78",x"08",x"00",x"17",x"42",x"01",x"00",x"07",x"71",x"d0",x"00",x"17",x"4f",x"40",x"10",x"ff",x"f9",x"91",x"00",x"08",x"00",x"0b",x"00",x"ba",x"f7",x"80",x"10",x"1a",x"04",x"00",x"0b",x"00",x"09",x"00",x"0e",x"00",x"eb",x"0a",x"00",x"89",x"24",x"78",x"08",x"00",x"13",x"07",x"00",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"20",x"17",x"42",x"00",x"08",x"31",x"00",x"09",x"00",x"98",x"07",x"40",x"10",x"31",x"21",x"40",x"10",x"4f",x"4f",x"10",x"4f",x"31",x"00",x"07",x"4f",x"5f",x"6f",x"72",x"14",x"24",x"07",x"7f",x"17",x"27",x"00",x"23",x"12",x"2c",x"14",x"ff",x"07",x"00",x"2f",x"f2",x"07",x"00",x"a0",x"10",x"ff",x"8f",x"18",x"0e",x"02",x"00",x"09",x"00",x"02",x"00",x"0a",x"00",x"a9",x"08",x"00",x"00",x"02",x"09",x"04",x"73",x"11",x"04",x"00",x"07",x"00",x"05",x"00",x"08",x"24",x"00",x"87",x"01",x"02",x"00",x"01",x"13",x"00",x"10",x"ef",x"1f",x"00",x"01",x"18",x"15",x"81",x"1c",x"0b",x"04",x"ea",x"41",x"01",x"4f",x"62",x"0d",x"02",x"64",x"02",x"4d",x"10",x"1f",x"01",x"54",x"06",x"62",x"0d",x"02",x"64",x"02",x"8d",x"10",x"1f",x"01",x"54",x"06",x"62",x"0d",x"02",x"64",x"02",x"cd",x"10",x"1f",x"01",x"21",x"ff",x"18",x"14",x"01",x"0c",x"4f",x"15",x"62",x"8d",x"10",x"03",x"05",x"21",x"32",x"15",x"cd",x"10",x"30",x"52",x"64",x"0c",x"2f",x"03",x"c2",x"e3",x"71",x"2f",x"5f",x"1f",x"6f",x"11",x"63",x"31",x"00",x"31",x"01",x"8d",x"10",x"34",x"52",x"cf",x"4d",x"10",x"34",x"02",x"c2",x"02",x"06",x"38",x"4d",x"10",x"01",x"61",x"34",x"2f",x"1c",x"01",x"0c",x"7f",x"61",x"33",x"71",x"01",x"15",x"1f",x"21",x"1f",x"2f",x"ff",x"f5",x"01",x"20",x"06",x"00",x"3f",x"32",x"3f",x"4f",x"0d",x"10",x"10",x"f6",x"22",x"12",x"10",x"ff",x"21",x"e3",x"e0",x"10",x"41",x"c0",x"10",x"01",x"52",x"31",x"55",x"12",x"2f",x"3f",x"4f",x"4d",x"10",x"10",x"c3",x"14",x"9f",x"ff",x"61",x"07",x"00",x"c0",x"10",x"1c",x"60",x"10",x"10",x"18",x"17",x"08",x"a3",x"40",x"10",x"b8",x"00",x"07",x"00",x"73",x"00",x"11",x"57",x"7f",x"73",x"02",x"0e",x"40",x"10",x"41",x"20",x"10",x"00",x"10",x"80",x"10",x"14",x"01",x"80",x"10",x"00",x"54",x"01",x"00",x"06",x"00",x"e0",x"10",x"80",x"10",x"01",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"18",x"00",x"00",x"01",x"19",x"10",x"01",x"80",x"10",x"a0",x"00",x"09",x"6f",x"5f",x"4f",x"df",x"ec",x"d0",x"e1",x"e1",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"02",x"18",x"06",x"f5",x"e2",x"f3",x"17",x"ce",x"06",x"10",x"00",x"60",x"10",x"10",x"10",x"c0",x"10",x"01",x"14",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"18",x"10",x"14",x"10",x"20",x"fb",x"41",x"7f",x"41",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"02",x"18",x"05",x"f5",x"42",x"f2",x"18",x"01",x"41",x"20",x"fa",x"4f",x"4f",x"5f",x"15",x"51",x"15",x"12",x"42",x"24",x"23",x"8d",x"10",x"02",x"04",x"08",x"22",x"21",x"01",x"d0",x"8f",x"4f",x"13",x"03",x"00",x"14",x"00",x"00",x"07",x"33",x"71",x"07",x"01",x"37",x"20",x"10",x"73",x"cd",x"10",x"10",x"07",x"00",x"73",x"cd",x"10",x"8d",x"10",x"4f",x"df",x"8f",x"10",x"13",x"f7",x"37",x"01",x"78",x"80",x"10",x"00",x"10",x"15",x"0b",x"04",x"00",x"02",x"03",x"31",x"31",x"10",x"8f",x"01",x"df",x"04",x"c0",x"10",x"01",x"13",x"31",x"04",x"13",x"31",x"10",x"f3",x"55",x"53",x"01",x"31",x"33",x"33",x"07",x"02",x"71",x"04",x"0f",x"f3",x"01",x"13",x"01",x"11",x"13",x"41",x"03",x"0d",x"10",x"00",x"c3",x"42",x"21",x"7f",x"4f",x"df",x"8f",x"10",x"07",x"07",x"00",x"32",x"21",x"01",x"10",x"a0",x"10",x"32",x"37",x"71",x"31",x"72",x"32",x"d0",x"4f",x"4f",x"5f",x"25",x"cd",x"10",x"01",x"04",x"01",x"08",x"cf",x"10",x"cf",x"4f",x"5f",x"6f",x"26",x"02",x"00",x"4b",x"37",x"2f",x"f2",x"27",x"20",x"14",x"ff",x"f2",x"08",x"7f",x"8f",x"2f",x"72",x"d2",x"80",x"10",x"20",x"e2",x"80",x"10",x"00",x"ff",x"f7",x"19",x"71",x"40",x"10",x"1a",x"ff",x"40",x"10",x"40",x"10",x"98",x"20",x"10",x"00",x"21",x"e0",x"10",x"04",x"17",x"40",x"10",x"18",x"ff",x"40",x"10",x"40",x"10",x"71",x"20",x"10",x"00",x"b6",x"a0",x"10",x"1f",x"b5",x"01",x"64",x"2c",x"52",x"04",x"1f",x"cf",x"62",x"03",x"18",x"0b",x"06",x"14",x"00",x"21",x"01",x"4f",x"8d",x"10",x"14",x"00",x"03",x"30",x"05",x"f8",x"21",x"01",x"11",x"30",x"4f",x"4d",x"10",x"2c",x"01",x"2f",x"21",x"1f",x"01",x"18",x"04",x"2f",x"7f",x"03",x"31",x"7f",x"31",x"72",x"02",x"31",x"00",x"01",x"07",x"28",x"12",x"20",x"24",x"3f",x"31",x"fc",x"00",x"11",x"10",x"ff",x"21",x"63",x"00",x"10",x"10",x"01",x"c0",x"10",x"10",x"07",x"1f",x"08",x"22",x"3f",x"6a",x"07",x"00",x"20",x"01",x"00",x"40",x"2f",x"ff",x"f2",x"14",x"21",x"01",x"3f",x"41",x"01",x"00",x"26",x"01",x"00",x"00",x"01",x"13",x"01",x"00",x"03",x"e0",x"10",x"9f",x"8f",x"17",x"11",x"1f",x"20",x"10",x"a0",x"10",x"14",x"01",x"80",x"10",x"01",x"4b",x"01",x"00",x"00",x"10",x"ff",x"f2",x"01",x"07",x"01",x"71",x"bf",x"71",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"15",x"40",x"10",x"53",x"a4",x"fc",x"02",x"20",x"cf",x"52",x"62",x"28",x"ec",x"c1",x"80",x"10",x"1f",x"4f",x"6f",x"3f",x"41",x"0d",x"10",x"20",x"21",x"20",x"24",x"14",x"21",x"1f",x"41",x"fb",x"af",x"c8",x"13",x"00",x"0a",x"00",x"07",x"14",x"40",x"10",x"40",x"10",x"7f",x"71",x"87",x"06",x"03",x"00",x"a1",x"01",x"00",x"11",x"61",x"23",x"10",x"40",x"06",x"6f",x"5f",x"4f",x"df",x"4f",x"10",x"01",x"1c",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"11",x"21",x"53",x"71",x"0d",x"10",x"1c",x"c1",x"51",x"ff",x"f4",x"00",x"60",x"8f",x"08",x"00",x"81",x"7f",x"81",x"02",x"12",x"21",x"08",x"12",x"21",x"21",x"aa",x"13",x"32",x"01",x"66",x"21",x"11",x"21",x"12",x"21",x"1e",x"21",x"02",x"12",x"14",x"a0",x"7f",x"5f",x"00",x"10",x"01",x"14",x"12",x"21",x"04",x"12",x"21",x"10",x"f2",x"55",x"52",x"01",x"21",x"33",x"32",x"03",x"02",x"31",x"04",x"0f",x"f2",x"01",x"12",x"01",x"11",x"21",x"43",x"81",x"8d",x"10",x"18",x"0c",x"41",x"1f",x"00",x"10",x"cf",x"10",x"10",x"01",x"89",x"17",x"00",x"14",x"12",x"4f",x"0e",x"09",x"10",x"32",x"8b",x"1e",x"29",x"91",x"88",x"21",x"98",x"11",x"87",x"71",x"d0",x"8f",x"00",x"df",x"04",x"8d",x"10",x"04",x"8f",x"10",x"03",x"20",x"10",x"a0",x"10",x"01",x"78",x"87",x"04",x"78",x"87",x"01",x"09",x"10",x"97",x"97",x"04",x"f7",x"0a",x"aa",x"ab",x"8b",x"0a",x"08",x"9b",x"9b",x"66",x"b7",x"0e",x"02",x"7b",x"b8",x"87",x"a7",x"a7",x"0a",x"02",x"a8",x"04",x"0f",x"f9",x"97",x"02",x"79",x"89",x"88",x"77",x"78",x"f8",x"00",x"60",x"10",x"10",x"07",x"03",x"08",x"03",x"00",x"81",x"07",x"ff",x"3b",x"aa",x"33",x"f8",x"ba",x"a1",x"bb",x"2b",x"9b",x"ea",x"40",x"10",x"01",x"03",x"d0",x"4f",x"4f",x"5f",x"25",x"cd",x"10",x"01",x"04",x"01",x"08",x"cf",x"10",x"b0",x"79",x"c1",x"99",x"d7",x"47",x"a4",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"74",x"63",x"61",x"74",x"00",x"70",x"6f",x"6e",x"72",x"70",x"6d",x"72",x"6f",x"6f",x"61",x"0a",x"20",x"69",x"69",x"72",x"70",x"6d",x"72",x"6f",x"6f",x"61",x"0a",x"6f",x"65",x"6e",x"74",x"20",x"20",x"61",x"65",x"66",x"63",x"6d",x"2e",x"4b",x"72",x"6d",x"65",x"6e",x"72",x"74",x"20",x"20",x"65",x"6b",x"32",x"61",x"61",x"6e",x"6e",x"72",x"74",x"20",x"20",x"65",x"6b",x"5b",x"45",x"52",x"69",x"63",x"30",x"34",x"20",x"75",x"62",x"78",x"78",x"25",x"52",x"21",x"74",x"20",x"20",x"30",x"2d",x"6f",x"20",x"30",x"34",x"5b",x"45",x"52",x"74",x"20",x"20",x"30",x"2d",x"6f",x"20",x"30",x"34",x"43",x"4d",x"20",x"65",x"20",x"6c",x"54",x"6c",x"63",x"20",x"20",x"6c",x"54",x"6c",x"6d",x"73",x"29",x"66",x"74",x"74",x"73",x"63",x"3a",x"0a",x"52",x"20",x"74",x"65",x"65",x"72",x"20",x"73",x"30",x"63",x"6f",x"20",x"69",x"65",x"74",x"49",x"61",x"6e",x"20",x"20",x"6c",x"43",x"69",x"20",x"73",x"20",x"73",x"43",x"32",x"43",x"61",x"6c",x"6c",x"20",x"20",x"67",x"45",x"53",x"33",x"6e",x"00",x"70",x"72",x"61",x"20",x"25",x"4d",x"72",x"6f",x"69",x"20",x"73",x"54",x"00",x"64",x"20",x"20",x"20",x"30",x"34",x"5b",x"63",x"69",x"20",x"20",x"30",x"34",x"5b",x"63",x"61",x"78",x"20",x"30",x"34",x"5b",x"63",x"74",x"20",x"20",x"30",x"34",x"5b",x"63",x"69",x"20",x"20",x"30",x"34",x"43",x"65",x"6f",x"61",x"6e",x"6c",x"74",x"20",x"20",x"64",x"74",x"66",x"72",x"61",x"72",x"72",x"67",x"6c",x"0a",x"72",x"72",x"2e",x"20",x"2f",x"20",x"20",x"73",x"72",x"20",x"65",x"64",x"61",x"74",x"6c",x"74",x"70",x"74",x"20",x"20",x"73",x"65",x"76",x"65",x"70",x"73",x"6f",x"72",x"69",x"72",x"6c",x"6f",x"20",x"77",x"6c",x"6f",x"0a",x"2e",x"31",x"54",x"2b",x"31",x"34",x"00",x"30",x"5e",x"35",x"2b",x"2e",x"65",x"2d",x"2b",x"00",x"36",x"32",x"2e",x"30",x"31",x"35",x"2d",x"2e",x"00",x"36",x"30",x"31",x"32",x"2d",x"00",x"32",x"55",x"00",x"33",x"37",x"62",x"66",x"6a",x"6e",x"72",x"76",x"7a",x"32",x"36",x"41",x"45",x"49",x"4d",x"51",x"55",x"59",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
 shared variable RAM3: RAM_TABLE := RAM_TABLE'(
x"81",x"70",x"ad",x"7e",x"70",x"90",x"10",x"70",x"81",x"70",x"40",x"ff",x"43",x"f6",x"89",x"80",x"70",x"70",x"50",x"10",x"cf",x"50",x"00",x"00",x"00",x"40",x"24",x"84",x"60",x"41",x"70",x"38",x"70",x"38",x"38",x"5e",x"90",x"90",x"90",x"90",x"0c",x"3a",x"40",x"60",x"42",x"77",x"ce",x"38",x"40",x"04",x"40",x"70",x"60",x"42",x"45",x"90",x"62",x"40",x"40",x"40",x"99",x"90",x"72",x"49",x"0c",x"3a",x"90",x"c8",x"38",x"99",x"80",x"60",x"41",x"91",x"44",x"60",x"42",x"42",x"90",x"80",x"99",x"ca",x"38",x"99",x"80",x"60",x"41",x"91",x"40",x"80",x"90",x"0c",x"80",x"7f",x"c2",x"38",x"80",x"70",x"40",x"40",x"77",x"05",x"98",x"11",x"40",x"40",x"40",x"52",x"38",x"5f",x"90",x"0c",x"40",x"90",x"0c",x"40",x"0c",x"0c",x"40",x"82",x"98",x"98",x"98",x"18",x"30",x"60",x"41",x"19",x"80",x"70",x"20",x"40",x"40",x"05",x"19",x"04",x"40",x"05",x"99",x"99",x"3a",x"82",x"30",x"19",x"99",x"91",x"30",x"5e",x"90",x"90",x"90",x"90",x"98",x"99",x"3a",x"60",x"40",x"44",x"c4",x"38",x"60",x"70",x"60",x"70",x"40",x"0c",x"40",x"90",x"70",x"40",x"3a",x"c0",x"38",x"38",x"40",x"20",x"40",x"c0",x"38",x"38",x"70",x"c3",x"38",x"38",x"20",x"98",x"9a",x"07",x"41",x"41",x"18",x"60",x"41",x"40",x"0c",x"38",x"70",x"c1",x"38",x"18",x"0c",x"cf",x"38",x"60",x"41",x"18",x"98",x"1a",x"40",x"00",x"40",x"38",x"40",x"3a",x"20",x"c1",x"38",x"40",x"40",x"04",x"90",x"18",x"60",x"42",x"18",x"18",x"10",x"60",x"50",x"89",x"06",x"3a",x"c0",x"38",x"40",x"40",x"90",x"98",x"40",x"70",x"70",x"90",x"88",x"60",x"20",x"45",x"98",x"0c",x"40",x"40",x"0c",x"40",x"18",x"98",x"90",x"98",x"90",x"90",x"18",x"10",x"10",x"c0",x"38",x"38",x"c5",x"38",x"60",x"04",x"98",x"99",x"07",x"42",x"18",x"ce",x"38",x"38",x"40",x"c1",x"38",x"98",x"9a",x"07",x"42",x"18",x"ce",x"38",x"60",x"42",x"80",x"7f",x"20",x"40",x"3a",x"40",x"18",x"60",x"41",x"98",x"18",x"40",x"40",x"40",x"40",x"18",x"10",x"ff",x"cf",x"38",x"18",x"c2",x"38",x"60",x"84",x"98",x"19",x"c3",x"38",x"0c",x"cd",x"38",x"60",x"98",x"98",x"04",x"40",x"52",x"38",x"99",x"3a",x"6f",x"43",x"43",x"60",x"42",x"80",x"7f",x"98",x"99",x"07",x"41",x"43",x"18",x"ce",x"38",x"38",x"c2",x"38",x"3a",x"40",x"40",x"c0",x"38",x"38",x"60",x"41",x"30",x"0c",x"38",x"30",x"70",x"c0",x"38",x"38",x"18",x"0c",x"cf",x"38",x"30",x"70",x"30",x"5d",x"70",x"90",x"90",x"90",x"90",x"90",x"90",x"60",x"41",x"c9",x"38",x"70",x"70",x"70",x"90",x"70",x"40",x"40",x"90",x"60",x"c1",x"38",x"40",x"0c",x"90",x"60",x"43",x"60",x"45",x"60",x"42",x"60",x"41",x"18",x"70",x"0c",x"38",x"c0",x"38",x"c4",x"38",x"5f",x"0c",x"40",x"c0",x"38",x"38",x"49",x"98",x"60",x"42",x"50",x"70",x"40",x"40",x"0c",x"46",x"45",x"90",x"0c",x"0c",x"40",x"40",x"40",x"40",x"38",x"c1",x"38",x"40",x"0c",x"0c",x"48",x"18",x"40",x"0c",x"5f",x"40",x"90",x"c2",x"38",x"40",x"40",x"70",x"50",x"c0",x"38",x"38",x"40",x"ce",x"38",x"40",x"38",x"40",x"90",x"0c",x"40",x"40",x"98",x"60",x"98",x"88",x"90",x"98",x"0c",x"43",x"98",x"98",x"98",x"18",x"30",x"cf",x"38",x"98",x"98",x"90",x"90",x"18",x"10",x"10",x"38",x"40",x"40",x"40",x"40",x"10",x"30",x"00",x"10",x"40",x"71",x"40",x"40",x"40",x"40",x"80",x"70",x"80",x"60",x"40",x"20",x"40",x"40",x"40",x"60",x"11",x"40",x"20",x"45",x"80",x"90",x"07",x"48",x"18",x"40",x"90",x"10",x"40",x"40",x"40",x"60",x"11",x"98",x"84",x"0c",x"38",x"90",x"c7",x"38",x"40",x"60",x"70",x"80",x"07",x"48",x"80",x"07",x"48",x"0c",x"77",x"20",x"20",x"40",x"85",x"88",x"85",x"18",x"10",x"40",x"90",x"0c",x"91",x"0c",x"40",x"07",x"49",x"18",x"60",x"42",x"98",x"98",x"80",x"7f",x"20",x"c9",x"38",x"f0",x"ff",x"80",x"07",x"49",x"88",x"06",x"04",x"98",x"91",x"18",x"60",x"cd",x"38",x"ff",x"70",x"40",x"98",x"98",x"98",x"18",x"30",x"5f",x"40",x"40",x"18",x"40",x"c3",x"38",x"98",x"50",x"c2",x"38",x"0c",x"10",x"18",x"40",x"50",x"98",x"19",x"99",x"91",x"98",x"0c",x"30",x"5f",x"90",x"0c",x"40",x"40",x"98",x"91",x"91",x"91",x"91",x"60",x"42",x"0c",x"c6",x"38",x"40",x"40",x"91",x"0c",x"c4",x"38",x"40",x"40",x"91",x"60",x"41",x"91",x"50",x"cb",x"38",x"40",x"40",x"40",x"70",x"30",x"00",x"40",x"90",x"90",x"90",x"90",x"8c",x"0c",x"40",x"60",x"40",x"80",x"90",x"c7",x"38",x"c9",x"38",x"40",x"c8",x"38",x"40",x"c8",x"38",x"40",x"c7",x"38",x"40",x"c6",x"38",x"60",x"42",x"0c",x"40",x"40",x"c0",x"38",x"38",x"40",x"60",x"41",x"99",x"70",x"c5",x"38",x"40",x"f1",x"91",x"91",x"91",x"43",x"60",x"41",x"99",x"70",x"c1",x"38",x"40",x"c1",x"38",x"76",x"40",x"40",x"40",x"40",x"40",x"80",x"90",x"90",x"91",x"91",x"70",x"84",x"70",x"04",x"60",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"60",x"40",x"00",x"60",x"04",x"40",x"40",x"80",x"98",x"0c",x"40",x"c0",x"38",x"90",x"80",x"98",x"60",x"42",x"70",x"20",x"04",x"90",x"80",x"98",x"80",x"98",x"60",x"42",x"80",x"7f",x"8b",x"00",x"40",x"c1",x"38",x"40",x"ca",x"38",x"40",x"40",x"04",x"c3",x"38",x"40",x"40",x"40",x"85",x"80",x"98",x"98",x"80",x"98",x"c5",x"38",x"40",x"04",x"c1",x"38",x"40",x"40",x"98",x"c6",x"38",x"40",x"cc",x"38",x"90",x"70",x"38",x"40",x"8b",x"90",x"c0",x"38",x"40",x"40",x"c0",x"38",x"40",x"c0",x"38",x"f0",x"70",x"80",x"90",x"0c",x"40",x"70",x"c0",x"38",x"80",x"98",x"0c",x"60",x"70",x"40",x"6f",x"c0",x"38",x"05",x"04",x"c0",x"38",x"40",x"80",x"98",x"0c",x"40",x"70",x"c0",x"38",x"70",x"40",x"98",x"50",x"20",x"40",x"40",x"8c",x"80",x"90",x"c4",x"38",x"40",x"c4",x"38",x"99",x"70",x"c9",x"38",x"99",x"3a",x"40",x"0c",x"40",x"c7",x"38",x"99",x"3a",x"40",x"0c",x"60",x"7f",x"40",x"47",x"ef",x"c0",x"38",x"38",x"40",x"40",x"70",x"38",x"40",x"42",x"80",x"6f",x"42",x"43",x"fe",x"c8",x"38",x"44",x"ea",x"cb",x"38",x"40",x"40",x"70",x"38",x"40",x"40",x"70",x"38",x"60",x"c9",x"38",x"40",x"40",x"70",x"40",x"18",x"c7",x"38",x"60",x"40",x"60",x"40",x"40",x"60",x"40",x"40",x"70",x"80",x"90",x"ff",x"00",x"60",x"40",x"40",x"70",x"60",x"40",x"60",x"40",x"60",x"40",x"80",x"98",x"8b",x"80",x"70",x"40",x"98",x"04",x"c0",x"38",x"43",x"99",x"80",x"98",x"19",x"07",x"42",x"f4",x"0c",x"40",x"99",x"50",x"40",x"40",x"04",x"c3",x"38",x"40",x"60",x"40",x"07",x"42",x"f7",x"0c",x"40",x"99",x"50",x"40",x"40",x"04",x"c2",x"38",x"40",x"60",x"40",x"07",x"42",x"fa",x"0c",x"40",x"99",x"50",x"40",x"60",x"40",x"60",x"40",x"50",x"60",x"84",x"f6",x"18",x"cf",x"38",x"60",x"40",x"60",x"40",x"60",x"40",x"60",x"40",x"60",x"40",x"60",x"40",x"60",x"40",x"40",x"80",x"90",x"fd",x"98",x"c7",x"38",x"40",x"c7",x"38",x"ca",x"38",x"f0",x"0c",x"40",x"0c",x"40",x"0c",x"70",x"80",x"90",x"c7",x"38",x"60",x"41",x"70",x"60",x"40",x"70",x"c5",x"38",x"70",x"45",x"70",x"80",x"98",x"70",x"60",x"41",x"f6",x"98",x"18",x"20",x"40",x"0c",x"0c",x"40",x"0c",x"0c",x"c7",x"38",x"f1",x"0c",x"40",x"0c",x"40",x"0c",x"60",x"70",x"80",x"90",x"cd",x"38",x"60",x"41",x"70",x"60",x"40",x"a4",x"70",x"cb",x"38",x"70",x"43",x"70",x"60",x"40",x"60",x"40",x"60",x"40",x"80",x"70",x"60",x"41",x"f3",x"c3",x"38",x"f6",x"98",x"18",x"20",x"40",x"40",x"f8",x"fa",x"c1",x"38",x"40",x"40",x"40",x"fe",x"f0",x"cf",x"38",x"40",x"ce",x"38",x"40",x"04",x"c0",x"38",x"60",x"40",x"38",x"60",x"40",x"60",x"42",x"80",x"98",x"70",x"40",x"74",x"20",x"99",x"f2",x"c9",x"38",x"80",x"7f",x"20",x"07",x"49",x"98",x"f6",x"70",x"60",x"42",x"18",x"c4",x"38",x"60",x"40",x"f6",x"70",x"8b",x"00",x"40",x"40",x"40",x"50",x"60",x"84",x"18",x"cd",x"38",x"40",x"04",x"40",x"18",x"60",x"40",x"42",x"60",x"42",x"70",x"40",x"74",x"8b",x"00",x"40",x"40",x"40",x"50",x"60",x"0c",x"20",x"07",x"49",x"60",x"42",x"70",x"40",x"74",x"8b",x"00",x"40",x"40",x"40",x"50",x"60",x"0c",x"20",x"07",x"49",x"80",x"98",x"80",x"7f",x"60",x"41",x"41",x"3a",x"c8",x"38",x"40",x"40",x"f9",x"c4",x"38",x"60",x"40",x"c7",x"38",x"40",x"40",x"8b",x"c6",x"38",x"80",x"98",x"0c",x"40",x"0c",x"0c",x"cb",x"38",x"f7",x"0c",x"40",x"40",x"40",x"40",x"ff",x"f0",x"ce",x"38",x"40",x"38",x"40",x"40",x"80",x"98",x"c2",x"38",x"40",x"40",x"40",x"70",x"40",x"38",x"5f",x"90",x"90",x"0c",x"40",x"40",x"40",x"90",x"0c",x"38",x"c0",x"38",x"40",x"40",x"51",x"38",x"98",x"10",x"40",x"40",x"0c",x"40",x"c5",x"38",x"40",x"90",x"70",x"20",x"80",x"50",x"88",x"00",x"00",x"ce",x"38",x"07",x"49",x"70",x"20",x"80",x"50",x"88",x"88",x"00",x"19",x"8b",x"10",x"49",x"50",x"cc",x"38",x"40",x"70",x"70",x"20",x"80",x"88",x"00",x"98",x"00",x"c0",x"38",x"70",x"38",x"07",x"43",x"70",x"50",x"07",x"49",x"50",x"07",x"49",x"3a",x"0c",x"40",x"98",x"0c",x"0c",x"40",x"20",x"70",x"10",x"20",x"40",x"07",x"40",x"00",x"19",x"3a",x"20",x"cd",x"38",x"10",x"cb",x"38",x"70",x"70",x"20",x"80",x"88",x"00",x"98",x"00",x"c0",x"38",x"70",x"38",x"70",x"c0",x"38",x"00",x"50",x"07",x"49",x"50",x"07",x"49",x"3a",x"c5",x"38",x"60",x"42",x"90",x"70",x"98",x"8b",x"70",x"20",x"70",x"88",x"00",x"8b",x"80",x"50",x"00",x"40",x"40",x"00",x"19",x"3a",x"20",x"cd",x"38",x"0c",x"07",x"49",x"50",x"ca",x"38",x"40",x"70",x"70",x"20",x"80",x"88",x"00",x"00",x"c0",x"38",x"70",x"38",x"70",x"c0",x"38",x"00",x"50",x"07",x"49",x"50",x"07",x"49",x"98",x"3a",x"c7",x"38",x"60",x"42",x"0c",x"40",x"77",x"90",x"98",x"8b",x"70",x"40",x"20",x"88",x"80",x"70",x"80",x"88",x"00",x"3a",x"20",x"07",x"88",x"00",x"3a",x"20",x"40",x"40",x"04",x"20",x"cc",x"38",x"50",x"40",x"ca",x"38",x"40",x"07",x"49",x"70",x"70",x"8b",x"70",x"20",x"40",x"18",x"40",x"07",x"46",x"50",x"41",x"70",x"c0",x"38",x"00",x"0c",x"cc",x"38",x"0c",x"cb",x"38",x"40",x"38",x"70",x"40",x"40",x"0c",x"c7",x"38",x"70",x"c6",x"38",x"3a",x"40",x"60",x"42",x"98",x"98",x"70",x"20",x"80",x"50",x"88",x"00",x"82",x"11",x"49",x"50",x"cd",x"38",x"38",x"c1",x"38",x"40",x"40",x"40",x"3a",x"30",x"60",x"42",x"70",x"20",x"80",x"50",x"88",x"00",x"00",x"ce",x"38",x"07",x"49",x"30",x"00",x"10",x"c3",x"38",x"8b",x"70",x"20",x"07",x"40",x"40",x"00",x"3a",x"20",x"cd",x"38",x"07",x"49",x"18",x"30",x"5f",x"90",x"10",x"c5",x"38",x"70",x"70",x"20",x"80",x"88",x"00",x"00",x"c0",x"38",x"70",x"38",x"07",x"43",x"70",x"50",x"07",x"49",x"50",x"07",x"49",x"18",x"40",x"50",x"38",x"90",x"10",x"c4",x"38",x"88",x"8b",x"70",x"00",x"80",x"88",x"50",x"88",x"00",x"19",x"3a",x"8b",x"00",x"49",x"50",x"07",x"49",x"18",x"40",x"30",x"5f",x"40",x"40",x"60",x"42",x"70",x"20",x"80",x"70",x"88",x"00",x"8b",x"80",x"50",x"00",x"40",x"40",x"00",x"19",x"3a",x"20",x"cd",x"38",x"10",x"cb",x"38",x"07",x"49",x"18",x"40",x"40",x"30",x"5e",x"40",x"40",x"90",x"60",x"42",x"70",x"70",x"20",x"90",x"98",x"80",x"70",x"88",x"80",x"10",x"20",x"20",x"07",x"88",x"88",x"00",x"19",x"3a",x"8b",x"89",x"89",x"04",x"8b",x"00",x"49",x"50",x"07",x"49",x"98",x"50",x"c8",x"38",x"98",x"98",x"51",x"38",x"5f",x"70",x"40",x"40",x"90",x"60",x"42",x"0c",x"60",x"42",x"70",x"80",x"8b",x"88",x"07",x"49",x"50",x"60",x"8b",x"c6",x"38",x"70",x"20",x"0c",x"20",x"70",x"8a",x"89",x"00",x"82",x"80",x"50",x"80",x"88",x"88",x"00",x"20",x"20",x"00",x"40",x"04",x"cb",x"38",x"00",x"ca",x"38",x"40",x"40",x"40",x"90",x"00",x"40",x"40",x"18",x"40",x"40",x"30",x"5a",x"90",x"90",x"0c",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"0c",x"40",x"60",x"41",x"43",x"8c",x"8c",x"ca",x"38",x"40",x"40",x"18",x"10",x"40",x"60",x"42",x"4d",x"98",x"0c",x"40",x"80",x"90",x"c2",x"38",x"1a",x"c0",x"38",x"12",x"07",x"49",x"90",x"90",x"0c",x"60",x"41",x"43",x"8c",x"8c",x"c2",x"38",x"40",x"40",x"18",x"10",x"40",x"60",x"42",x"4d",x"90",x"98",x"60",x"45",x"98",x"1a",x"c0",x"38",x"12",x"07",x"49",x"90",x"98",x"98",x"ce",x"38",x"98",x"cd",x"38",x"98",x"cc",x"38",x"98",x"cc",x"38",x"98",x"cb",x"38",x"98",x"ca",x"38",x"98",x"c9",x"38",x"98",x"c9",x"38",x"98",x"c8",x"38",x"98",x"c7",x"38",x"98",x"c6",x"38",x"98",x"c6",x"38",x"98",x"c5",x"38",x"98",x"c4",x"38",x"98",x"c3",x"38",x"98",x"c3",x"38",x"40",x"40",x"40",x"55",x"38",x"18",x"1a",x"c0",x"38",x"40",x"70",x"40",x"84",x"62",x"41",x"cc",x"38",x"c3",x"38",x"c9",x"38",x"c0",x"38",x"40",x"80",x"04",x"c1",x"38",x"40",x"90",x"70",x"40",x"60",x"47",x"60",x"42",x"ca",x"38",x"c0",x"38",x"40",x"90",x"70",x"40",x"60",x"42",x"ca",x"38",x"40",x"90",x"80",x"84",x"70",x"c0",x"38",x"40",x"80",x"84",x"70",x"ce",x"38",x"62",x"42",x"62",x"42",x"62",x"41",x"70",x"40",x"60",x"41",x"62",x"42",x"62",x"41",x"98",x"50",x"40",x"ca",x"38",x"c9",x"38",x"20",x"66",x"41",x"98",x"50",x"40",x"47",x"60",x"41",x"80",x"84",x"70",x"c6",x"38",x"40",x"98",x"62",x"90",x"70",x"42",x"70",x"38",x"40",x"20",x"60",x"49",x"47",x"80",x"84",x"70",x"c1",x"38",x"38",x"40",x"90",x"70",x"50",x"9a",x"80",x"60",x"42",x"0c",x"c3",x"38",x"38",x"40",x"80",x"10",x"30",x"98",x"50",x"40",x"38",x"40",x"90",x"41",x"98",x"50",x"40",x"38",x"40",x"90",x"80",x"70",x"38",x"10",x"40",x"40",x"40",x"40",x"40",x"72",x"70",x"38",x"20",x"18",x"85",x"80",x"80",x"07",x"49",x"cb",x"38",x"60",x"42",x"80",x"80",x"50",x"00",x"12",x"49",x"00",x"20",x"50",x"3a",x"20",x"c1",x"38",x"c4",x"38",x"40",x"c9",x"38",x"38",x"40",x"c1",x"38",x"c8",x"38",x"40",x"04",x"40",x"40",x"89",x"70",x"f3",x"c5",x"38",x"40",x"04",x"40",x"20",x"18",x"40",x"89",x"70",x"f2",x"c2",x"38",x"40",x"c1",x"38",x"20",x"20",x"70",x"40",x"98",x"98",x"98",x"18",x"30",x"0c",x"60",x"47",x"60",x"42",x"42",x"fb",x"44",x"60",x"42",x"60",x"42",x"42",x"f5",x"42",x"60",x"41",x"fb",x"41",x"f5",x"40",x"60",x"41",x"fb",x"18",x"38",x"40",x"20",x"84",x"60",x"42",x"06",x"40",x"40",x"05",x"40",x"20",x"c0",x"38",x"80",x"7f",x"40",x"89",x"85",x"89",x"06",x"20",x"c0",x"38",x"04",x"40",x"40",x"20",x"40",x"84",x"60",x"42",x"06",x"88",x"89",x"85",x"89",x"06",x"20",x"c0",x"38",x"04",x"40",x"40",x"20",x"40",x"84",x"60",x"42",x"06",x"88",x"89",x"85",x"89",x"06",x"20",x"c0",x"38",x"04",x"40",x"40",x"84",x"88",x"60",x"c0",x"38",x"04",x"40",x"40",x"80",x"7f",x"30",x"5f",x"90",x"0c",x"40",x"cc",x"38",x"89",x"cc",x"38",x"40",x"50",x"38",x"10",x"40",x"40",x"ff",x"84",x"c9",x"38",x"80",x"70",x"89",x"c8",x"38",x"89",x"04",x"40",x"0c",x"40",x"40",x"98",x"98",x"18",x"30",x"5f",x"90",x"0c",x"40",x"c4",x"38",x"80",x"70",x"89",x"c3",x"38",x"40",x"50",x"38",x"30",x"70",x"40",x"60",x"41",x"10",x"38",x"40",x"18",x"40",x"60",x"41",x"10",x"38",x"40",x"90",x"90",x"90",x"80",x"90",x"80",x"90",x"80",x"90",x"82",x"0c",x"60",x"80",x"90",x"80",x"90",x"80",x"0c",x"60",x"40",x"80",x"90",x"40",x"80",x"1a",x"c6",x"38",x"70",x"40",x"70",x"38",x"0c",x"40",x"40",x"62",x"47",x"62",x"42",x"42",x"05",x"4d",x"62",x"42",x"63",x"42",x"41",x"05",x"4c",x"62",x"41",x"72",x"38",x"4a",x"62",x"41",x"71",x"38",x"40",x"04",x"c2",x"38",x"40",x"20",x"50",x"80",x"80",x"0c",x"60",x"49",x"44",x"7f",x"62",x"41",x"80",x"98",x"7f",x"04",x"40",x"60",x"40",x"80",x"6f",x"43",x"71",x"70",x"20",x"7f",x"c0",x"38",x"38",x"60",x"40",x"60",x"40",x"40",x"40",x"40",x"20",x"60",x"47",x"0c",x"40",x"20",x"50",x"80",x"80",x"0c",x"60",x"49",x"45",x"80",x"90",x"80",x"90",x"80",x"90",x"7f",x"38",x"84",x"62",x"41",x"80",x"98",x"7f",x"40",x"04",x"40",x"60",x"40",x"9a",x"70",x"60",x"40",x"c0",x"38",x"72",x"04",x"c0",x"38",x"38",x"60",x"40",x"40",x"80",x"90",x"38",x"38",x"38",x"66",x"47",x"66",x"47",x"64",x"42",x"65",x"42",x"cf",x"38",x"60",x"40",x"05",x"60",x"40",x"38",x"c4",x"38",x"c2",x"38",x"c0",x"38",x"40",x"70",x"38",x"c1",x"38",x"c0",x"38",x"40",x"80",x"98",x"70",x"80",x"90",x"42",x"67",x"42",x"67",x"42",x"67",x"42",x"cb",x"38",x"80",x"98",x"7f",x"04",x"40",x"60",x"40",x"80",x"98",x"90",x"90",x"0c",x"60",x"40",x"40",x"0c",x"60",x"40",x"40",x"80",x"98",x"74",x"80",x"90",x"41",x"66",x"42",x"c4",x"38",x"60",x"40",x"70",x"80",x"98",x"50",x"80",x"80",x"90",x"70",x"80",x"90",x"c0",x"38",x"40",x"80",x"98",x"80",x"98",x"74",x"40",x"60",x"42",x"f1",x"80",x"98",x"70",x"1a",x"20",x"40",x"00",x"1a",x"40",x"40",x"40",x"40",x"40",x"00",x"1a",x"40",x"92",x"92",x"9a",x"89",x"04",x"00",x"92",x"1a",x"40",x"40",x"40",x"40",x"00",x"1a",x"40",x"92",x"92",x"9a",x"89",x"04",x"00",x"92",x"1a",x"40",x"40",x"40",x"40",x"00",x"1a",x"40",x"92",x"71",x"60",x"40",x"60",x"42",x"c5",x"38",x"60",x"40",x"c0",x"38",x"40",x"5e",x"72",x"ca",x"38",x"40",x"71",x"40",x"60",x"41",x"0c",x"38",x"40",x"80",x"00",x"80",x"98",x"80",x"90",x"00",x"60",x"41",x"8c",x"73",x"cc",x"38",x"c5",x"38",x"40",x"80",x"90",x"80",x"0c",x"40",x"ff",x"76",x"1a",x"0c",x"40",x"70",x"c9",x"38",x"70",x"92",x"0c",x"40",x"80",x"98",x"0c",x"45",x"60",x"48",x"44",x"8c",x"70",x"60",x"40",x"20",x"c5",x"38",x"40",x"00",x"12",x"c6",x"38",x"60",x"40",x"50",x"38",x"40",x"40",x"40",x"00",x"1a",x"80",x"98",x"80",x"50",x"ce",x"38",x"60",x"40",x"04",x"c0",x"38",x"40",x"80",x"98",x"80",x"98",x"80",x"07",x"45",x"c4",x"38",x"20",x"72",x"60",x"40",x"c2",x"38",x"60",x"40",x"80",x"90",x"c1",x"38",x"c4",x"38",x"60",x"40",x"50",x"80",x"80",x"90",x"80",x"98",x"70",x"c0",x"38",x"80",x"98",x"70",x"18",x"40",x"40",x"42",x"80",x"98",x"0c",x"c1",x"38",x"c0",x"38",x"60",x"40",x"04",x"c0",x"38",x"40",x"80",x"98",x"80",x"98",x"80",x"60",x"44",x"c0",x"38",x"72",x"c5",x"38",x"60",x"40",x"50",x"80",x"80",x"90",x"80",x"00",x"12",x"40",x"66",x"41",x"80",x"98",x"7f",x"50",x"70",x"80",x"90",x"18",x"60",x"40",x"60",x"40",x"40",x"60",x"40",x"60",x"40",x"05",x"60",x"41",x"cb",x"38",x"80",x"90",x"04",x"40",x"72",x"62",x"41",x"80",x"98",x"cf",x"38",x"60",x"40",x"50",x"80",x"80",x"90",x"18",x"c0",x"38",x"40",x"0c",x"c2",x"38",x"0c",x"c1",x"38",x"40",x"40",x"c0",x"38",x"0c",x"ce",x"38",x"60",x"40",x"82",x"04",x"c3",x"38",x"60",x"40",x"c0",x"38",x"40",x"00",x"82",x"0c",x"60",x"40",x"60",x"40",x"40",x"80",x"98",x"7f",x"00",x"60",x"40",x"60",x"40",x"ce",x"38",x"12",x"80",x"98",x"1a",x"c0",x"38",x"38",x"40",x"c9",x"38",x"50",x"40",x"40",x"60",x"42",x"12",x"50",x"40",x"80",x"98",x"80",x"98",x"42",x"80",x"98",x"cc",x"38",x"60",x"40",x"40",x"0c",x"60",x"40",x"80",x"60",x"04",x"40",x"60",x"40",x"12",x"40",x"44",x"0c",x"40",x"40",x"80",x"90",x"88",x"80",x"90",x"70",x"80",x"90",x"18",x"60",x"40",x"60",x"40",x"40",x"70",x"c0",x"38",x"80",x"98",x"71",x"70",x"80",x"90",x"80",x"98",x"80",x"98",x"c6",x"38",x"70",x"43",x"70",x"60",x"40",x"05",x"80",x"90",x"70",x"80",x"98",x"60",x"80",x"98",x"70",x"41",x"80",x"98",x"80",x"70",x"ff",x"06",x"60",x"40",x"60",x"40",x"cc",x"38",x"ff",x"04",x"c0",x"38",x"40",x"88",x"72",x"40",x"84",x"80",x"98",x"89",x"82",x"c8",x"38",x"80",x"90",x"60",x"45",x"1a",x"0c",x"12",x"c1",x"38",x"40",x"50",x"40",x"07",x"45",x"00",x"60",x"40",x"07",x"44",x"82",x"80",x"c0",x"38",x"12",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"9a",x"92",x"80",x"c0",x"38",x"38",x"40",x"cc",x"38",x"80",x"ce",x"38",x"60",x"40",x"0c",x"c2",x"38",x"40",x"50",x"1a",x"50",x"45",x"0c",x"c0",x"38",x"00",x"60",x"40",x"07",x"44",x"7f",x"80",x"0c",x"0c",x"40",x"00",x"60",x"40",x"c7",x"38",x"60",x"40",x"5f",x"60",x"45",x"0c",x"60",x"40",x"70",x"04",x"0c",x"41",x"80",x"70",x"0c",x"60",x"40",x"60",x"40",x"60",x"40",x"c7",x"38",x"ff",x"66",x"60",x"40",x"42",x"80",x"98",x"66",x"41",x"8c",x"8c",x"90",x"8c",x"90",x"80",x"98",x"80",x"98",x"80",x"98",x"0c",x"40",x"98",x"0c",x"c0",x"38",x"c9",x"38",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"60",x"40",x"60",x"40",x"40",x"98",x"60",x"41",x"80",x"0c",x"38",x"80",x"92",x"80",x"98",x"1a",x"12",x"60",x"40",x"44",x"41",x"72",x"40",x"40",x"38",x"40",x"c2",x"38",x"60",x"40",x"00",x"1a",x"12",x"07",x"41",x"74",x"c0",x"38",x"80",x"80",x"90",x"12",x"40",x"c2",x"38",x"60",x"40",x"60",x"40",x"70",x"40",x"7f",x"c0",x"38",x"40",x"80",x"70",x"40",x"80",x"90",x"c1",x"38",x"60",x"40",x"82",x"00",x"41",x"80",x"98",x"72",x"12",x"70",x"40",x"80",x"98",x"53",x"92",x"0c",x"40",x"70",x"40",x"53",x"92",x"80",x"98",x"00",x"ce",x"38",x"cd",x"38",x"80",x"ff",x"12",x"72",x"80",x"98",x"80",x"98",x"04",x"60",x"40",x"c9",x"38",x"80",x"98",x"c8",x"38",x"38",x"1a",x"c1",x"38",x"c6",x"38",x"c6",x"38",x"38",x"40",x"c0",x"38",x"cc",x"38",x"80",x"9a",x"60",x"42",x"5f",x"60",x"41",x"82",x"60",x"45",x"80",x"5f",x"1a",x"40",x"43",x"40",x"92",x"72",x"84",x"66",x"41",x"60",x"41",x"70",x"60",x"70",x"70",x"c0",x"38",x"50",x"62",x"42",x"04",x"cd",x"38",x"60",x"42",x"40",x"50",x"1a",x"c1",x"38",x"c0",x"38",x"ce",x"38",x"0c",x"40",x"40",x"cf",x"38",x"c0",x"38",x"40",x"c1",x"38",x"80",x"0c",x"20",x"20",x"40",x"ca",x"38",x"60",x"40",x"60",x"40",x"60",x"40",x"60",x"f0",x"0c",x"0c",x"42",x"80",x"9a",x"60",x"42",x"5f",x"60",x"41",x"82",x"71",x"20",x"60",x"41",x"60",x"44",x"43",x"80",x"0c",x"60",x"40",x"82",x"72",x"0c",x"40",x"80",x"98",x"00",x"80",x"90",x"40",x"5f",x"60",x"40",x"40",x"60",x"42",x"80",x"98",x"12",x"80",x"90",x"71",x"60",x"41",x"60",x"44",x"43",x"80",x"98",x"80",x"98",x"ff",x"0c",x"0c",x"40",x"00",x"80",x"90",x"40",x"5f",x"60",x"40",x"60",x"40",x"60",x"43",x"80",x"98",x"42",x"50",x"60",x"00",x"07",x"12",x"44",x"4e",x"80",x"98",x"00",x"60",x"45",x"0c",x"0c",x"40",x"00",x"40",x"40",x"82",x"8c",x"8c",x"0c",x"40",x"40",x"40",x"60",x"40",x"60",x"40",x"40",x"98",x"60",x"41",x"80",x"0c",x"38",x"80",x"92",x"80",x"98",x"1a",x"c0",x"38",x"38",x"60",x"c0",x"38",x"40",x"72",x"0c",x"40",x"40",x"40",x"80",x"80",x"c7",x"38",x"40",x"60",x"43",x"72",x"60",x"92",x"12",x"70",x"45",x"41",x"12",x"50",x"40",x"20",x"ce",x"38",x"60",x"42",x"12",x"40",x"9a",x"0c",x"c1",x"38",x"38",x"40",x"50",x"c0",x"38",x"12",x"1a",x"50",x"40",x"ce",x"38",x"38",x"cd",x"38",x"12",x"60",x"40",x"c3",x"38",x"60",x"f5",x"70",x"98",x"04",x"cf",x"38",x"50",x"80",x"9a",x"0c",x"cd",x"38",x"40",x"40",x"40",x"d1",x"30",x"00",x"10",x"40",x"40",x"40",x"0c",x"98",x"0c",x"60",x"42",x"7f",x"20",x"ff",x"04",x"c0",x"38",x"40",x"80",x"62",x"47",x"70",x"04",x"c4",x"38",x"c0",x"38",x"38",x"04",x"c1",x"38",x"72",x"38",x"5f",x"82",x"41",x"88",x"72",x"40",x"70",x"89",x"82",x"72",x"40",x"20",x"90",x"c0",x"38",x"38",x"c0",x"38",x"38",x"90",x"41",x"90",x"41",x"90",x"61",x"41",x"5f",x"88",x"71",x"40",x"40",x"04",x"90",x"c4",x"38",x"0c",x"40",x"40",x"0c",x"90",x"0c",x"40",x"98",x"00",x"98",x"12",x"0c",x"40",x"0c",x"60",x"41",x"40",x"73",x"0c",x"40",x"40",x"98",x"07",x"43",x"0c",x"40",x"40",x"40",x"40",x"20",x"04",x"c2",x"38",x"c0",x"38",x"38",x"72",x"cf",x"38",x"7f",x"38",x"98",x"ff",x"04",x"c0",x"38",x"50",x"40",x"60",x"42",x"61",x"42",x"41",x"77",x"40",x"12",x"41",x"60",x"41",x"73",x"50",x"40",x"40",x"04",x"c2",x"38",x"c0",x"38",x"38",x"40",x"40",x"0c",x"0c",x"40",x"00",x"40",x"5f",x"40",x"c2",x"38",x"82",x"73",x"0c",x"c3",x"38",x"98",x"00",x"60",x"46",x"0c",x"5f",x"40",x"00",x"12",x"ce",x"38",x"60",x"44",x"41",x"0c",x"0c",x"cf",x"38",x"20",x"38",x"98",x"98",x"98",x"18",x"30",x"5e",x"10",x"40",x"40",x"40",x"40",x"40",x"40",x"38",x"40",x"51",x"38",x"10",x"40",x"40",x"40",x"40",x"70",x"90",x"90",x"c4",x"38",x"60",x"41",x"70",x"40",x"40",x"70",x"40",x"6f",x"c0",x"38",x"98",x"05",x"60",x"45",x"0c",x"64",x"20",x"40",x"c0",x"38",x"90",x"98",x"60",x"c0",x"38",x"10",x"70",x"06",x"40",x"40",x"40",x"90",x"90",x"70",x"70",x"40",x"40",x"40",x"40",x"40",x"60",x"42",x"98",x"70",x"40",x"40",x"40",x"40",x"40",x"60",x"70",x"40",x"8c",x"0c",x"40",x"0c",x"60",x"85",x"7b",x"40",x"40",x"40",x"0c",x"60",x"70",x"40",x"0c",x"40",x"53",x"70",x"40",x"40",x"40",x"40",x"40",x"40",x"98",x"98",x"60",x"40",x"50",x"41",x"98",x"07",x"49",x"ce",x"38",x"40",x"1a",x"12",x"07",x"49",x"98",x"98",x"cd",x"38",x"40",x"40",x"70",x"40",x"60",x"c0",x"38",x"90",x"70",x"98",x"98",x"c8",x"38",x"70",x"45",x"70",x"40",x"70",x"60",x"42",x"47",x"98",x"98",x"a4",x"70",x"90",x"90",x"90",x"c6",x"38",x"f0",x"70",x"90",x"0c",x"40",x"98",x"60",x"40",x"80",x"cb",x"38",x"40",x"40",x"40",x"40",x"40",x"41",x"98",x"98",x"40",x"98",x"98",x"70",x"40",x"0c",x"40",x"40",x"60",x"42",x"70",x"40",x"60",x"45",x"80",x"90",x"07",x"40",x"47",x"98",x"55",x"90",x"c5",x"38",x"40",x"a4",x"70",x"0c",x"40",x"8c",x"0c",x"40",x"90",x"0c",x"40",x"40",x"40",x"98",x"53",x"12",x"07",x"47",x"98",x"07",x"49",x"98",x"65",x"45",x"42",x"1a",x"40",x"73",x"0c",x"12",x"40",x"38",x"12",x"38",x"40",x"92",x"44",x"9a",x"50",x"40",x"1a",x"63",x"45",x"12",x"c0",x"38",x"38",x"60",x"50",x"cd",x"38",x"c0",x"38",x"50",x"38",x"12",x"40",x"40",x"40",x"53",x"38",x"5e",x"10",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"98",x"18",x"30",x"00",x"f6",x"10",x"40",x"40",x"40",x"40",x"40",x"40",x"98",x"18",x"30",x"00",x"98",x"10",x"40",x"40",x"40",x"40",x"40",x"40",x"98",x"18",x"30",x"30",x"30",x"30",x"70",x"38",x"5f",x"90",x"cf",x"38",x"96",x"76",x"c5",x"38",x"40",x"50",x"38",x"70",x"30",x"70",x"30",x"70",x"20",x"c0",x"38",x"38",x"60",x"42",x"12",x"5f",x"20",x"ce",x"38",x"38",x"60",x"49",x"ff",x"60",x"88",x"05",x"40",x"c2",x"38",x"90",x"90",x"90",x"5f",x"60",x"47",x"40",x"10",x"5f",x"cf",x"38",x"c1",x"38",x"5f",x"60",x"41",x"30",x"5f",x"40",x"40",x"90",x"04",x"70",x"61",x"43",x"6f",x"43",x"c8",x"38",x"60",x"89",x"84",x"05",x"c0",x"38",x"38",x"70",x"04",x"90",x"0c",x"38",x"c3",x"38",x"70",x"7f",x"20",x"20",x"c1",x"38",x"10",x"20",x"40",x"c3",x"38",x"42",x"10",x"40",x"70",x"04",x"41",x"80",x"70",x"10",x"40",x"40",x"0c",x"30",x"5d",x"90",x"90",x"0c",x"0c",x"60",x"90",x"8e",x"84",x"81",x"70",x"60",x"70",x"47",x"70",x"70",x"42",x"70",x"42",x"0c",x"20",x"20",x"c3",x"38",x"8e",x"81",x"70",x"60",x"70",x"49",x"70",x"70",x"41",x"70",x"42",x"0c",x"60",x"41",x"70",x"60",x"42",x"70",x"f0",x"60",x"49",x"70",x"42",x"0c",x"60",x"41",x"88",x"70",x"05",x"c3",x"38",x"70",x"c0",x"38",x"70",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c1",x"38",x"60",x"0c",x"0c",x"40",x"f0",x"70",x"20",x"60",x"41",x"86",x"80",x"70",x"20",x"05",x"60",x"60",x"42",x"0c",x"c0",x"38",x"0c",x"40",x"06",x"60",x"41",x"0c",x"0c",x"40",x"85",x"60",x"41",x"c2",x"38",x"20",x"60",x"c6",x"38",x"70",x"c0",x"38",x"07",x"47",x"70",x"42",x"0c",x"60",x"41",x"0c",x"41",x"0c",x"c0",x"38",x"c0",x"38",x"ff",x"89",x"0c",x"20",x"60",x"60",x"20",x"42",x"90",x"cf",x"38",x"40",x"c6",x"38",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"40",x"38",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"89",x"85",x"80",x"0c",x"c2",x"38",x"70",x"82",x"89",x"ff",x"90",x"84",x"8f",x"7f",x"04",x"42",x"90",x"90",x"cf",x"38",x"40",x"c6",x"38",x"40",x"40",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"89",x"46",x"89",x"0c",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"89",x"85",x"80",x"0c",x"40",x"70",x"0c",x"20",x"40",x"40",x"40",x"05",x"60",x"85",x"c0",x"38",x"0c",x"38",x"20",x"70",x"c4",x"38",x"0c",x"40",x"40",x"40",x"90",x"0c",x"98",x"82",x"0c",x"40",x"85",x"70",x"c0",x"38",x"98",x"98",x"05",x"40",x"40",x"20",x"70",x"6f",x"90",x"98",x"98",x"88",x"89",x"05",x"40",x"60",x"05",x"43",x"43",x"8e",x"81",x"80",x"70",x"60",x"42",x"88",x"89",x"00",x"89",x"50",x"04",x"20",x"40",x"0c",x"06",x"0f",x"85",x"70",x"60",x"42",x"ff",x"6f",x"47",x"90",x"60",x"42",x"89",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"89",x"c8",x"38",x"20",x"60",x"c4",x"38",x"20",x"20",x"c3",x"38",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"89",x"05",x"40",x"0c",x"cd",x"38",x"40",x"0c",x"20",x"40",x"45",x"98",x"f0",x"70",x"0c",x"c9",x"38",x"c3",x"38",x"74",x"20",x"20",x"90",x"0c",x"40",x"05",x"c0",x"38",x"98",x"0c",x"c6",x"38",x"85",x"70",x"40",x"60",x"89",x"70",x"04",x"40",x"70",x"98",x"05",x"40",x"70",x"60",x"47",x"70",x"81",x"60",x"41",x"70",x"04",x"01",x"98",x"98",x"98",x"18",x"30",x"72",x"60",x"42",x"80",x"70",x"20",x"42",x"60",x"42",x"72",x"20",x"20",x"20",x"20",x"05",x"0c",x"38",x"5f",x"70",x"60",x"41",x"70",x"60",x"70",x"20",x"60",x"c0",x"38",x"c0",x"38",x"04",x"cb",x"38",x"70",x"60",x"41",x"70",x"f0",x"60",x"47",x"70",x"42",x"0c",x"60",x"41",x"85",x"85",x"05",x"60",x"42",x"84",x"60",x"45",x"70",x"07",x"49",x"70",x"07",x"45",x"70",x"42",x"42",x"70",x"07",x"47",x"70",x"07",x"43",x"70",x"42",x"0c",x"7f",x"c1",x"38",x"06",x"05",x"c0",x"38",x"18",x"50",x"38",x"5f",x"70",x"60",x"41",x"70",x"60",x"70",x"20",x"60",x"c0",x"38",x"c0",x"38",x"04",x"60",x"41",x"04",x"70",x"c0",x"38",x"70",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c8",x"38",x"20",x"20",x"70",x"c7",x"38",x"20",x"c2",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c2",x"38",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c0",x"38",x"04",x"7f",x"41",x"70",x"06",x"60",x"41",x"70",x"0c",x"30",x"5f",x"60",x"60",x"10",x"70",x"41",x"70",x"60",x"70",x"47",x"70",x"42",x"0c",x"60",x"41",x"ff",x"7f",x"60",x"70",x"41",x"70",x"60",x"c0",x"38",x"c0",x"38",x"18",x"30",x"00",x"70",x"10",x"c0",x"38",x"ff",x"7f",x"84",x"f0",x"60",x"47",x"70",x"42",x"0c",x"60",x"41",x"04",x"70",x"c0",x"38",x"70",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c8",x"38",x"20",x"20",x"70",x"c7",x"38",x"20",x"c2",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c2",x"38",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c0",x"38",x"04",x"60",x"41",x"70",x"06",x"60",x"41",x"70",x"0c",x"30",x"00",x"70",x"10",x"c0",x"38",x"ff",x"7f",x"84",x"f0",x"60",x"47",x"70",x"42",x"0c",x"60",x"41",x"04",x"70",x"c0",x"38",x"70",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c8",x"38",x"20",x"20",x"70",x"c7",x"38",x"20",x"c2",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c2",x"38",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c0",x"38",x"04",x"60",x"41",x"70",x"06",x"60",x"41",x"70",x"0c",x"30",x"00",x"70",x"10",x"c0",x"38",x"ff",x"7f",x"84",x"f0",x"60",x"47",x"70",x"42",x"0c",x"60",x"41",x"04",x"70",x"c0",x"38",x"70",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c8",x"38",x"20",x"20",x"70",x"c7",x"38",x"20",x"c2",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c2",x"38",x"38",x"70",x"c0",x"38",x"70",x"c0",x"38",x"c0",x"38",x"04",x"60",x"41",x"70",x"06",x"60",x"41",x"70",x"0c",x"30",x"00",x"70",x"10",x"c0",x"38",x"ff",x"7f",x"84",x"f0",x"60",x"47",x"70",x"42",x"0c",x"7f",x"cb",x"38",x"70",x"60",x"41",x"70",x"f0",x"60",x"47",x"70",x"42",x"0c",x"60",x"41",x"85",x"85",x"05",x"60",x"42",x"84",x"60",x"45",x"70",x"07",x"49",x"70",x"07",x"45",x"70",x"42",x"42",x"70",x"07",x"47",x"70",x"07",x"43",x"70",x"42",x"0c",x"60",x"c1",x"38",x"06",x"05",x"c0",x"38",x"18",x"50",x"38",x"5c",x"86",x"80",x"70",x"90",x"90",x"90",x"04",x"40",x"40",x"40",x"90",x"89",x"04",x"60",x"84",x"04",x"40",x"40",x"40",x"40",x"47",x"98",x"5f",x"40",x"48",x"c9",x"38",x"60",x"90",x"70",x"60",x"20",x"42",x"70",x"f0",x"60",x"49",x"70",x"42",x"0c",x"60",x"41",x"88",x"70",x"20",x"40",x"84",x"70",x"60",x"42",x"70",x"f0",x"60",x"49",x"70",x"40",x"42",x"0c",x"60",x"41",x"88",x"70",x"85",x"cc",x"38",x"90",x"90",x"90",x"70",x"40",x"40",x"05",x"40",x"40",x"20",x"60",x"82",x"70",x"90",x"0c",x"40",x"70",x"0c",x"20",x"c7",x"38",x"40",x"40",x"0c",x"20",x"0c",x"40",x"70",x"0c",x"20",x"c4",x"38",x"40",x"40",x"0c",x"20",x"0c",x"40",x"70",x"0c",x"20",x"c1",x"38",x"40",x"40",x"05",x"40",x"40",x"88",x"70",x"40",x"98",x"0c",x"0c",x"ce",x"38",x"20",x"70",x"01",x"0f",x"03",x"cc",x"38",x"40",x"0c",x"0c",x"40",x"98",x"70",x"0e",x"7f",x"81",x"90",x"90",x"98",x"98",x"88",x"89",x"05",x"60",x"85",x"70",x"c7",x"38",x"40",x"0c",x"90",x"c6",x"38",x"40",x"40",x"8e",x"70",x"20",x"40",x"c4",x"38",x"70",x"01",x"40",x"98",x"84",x"70",x"40",x"98",x"0e",x"81",x"0e",x"20",x"8e",x"98",x"81",x"98",x"98",x"9f",x"6f",x"20",x"40",x"20",x"47",x"90",x"0c",x"98",x"98",x"cd",x"38",x"40",x"5f",x"88",x"03",x"38",x"60",x"86",x"05",x"cb",x"38",x"05",x"c6",x"38",x"40",x"88",x"89",x"89",x"05",x"90",x"98",x"98",x"c7",x"38",x"40",x"0f",x"40",x"98",x"83",x"00",x"40",x"45",x"c1",x"38",x"40",x"c0",x"38",x"38",x"40",x"70",x"20",x"07",x"c0",x"38",x"07",x"47",x"70",x"42",x"0c",x"60",x"88",x"04",x"98",x"0e",x"70",x"20",x"ce",x"38",x"05",x"c1",x"38",x"cd",x"38",x"cc",x"38",x"40",x"20",x"c0",x"38",x"40",x"85",x"60",x"42",x"70",x"60",x"c2",x"38",x"ca",x"38",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"40",x"40",x"f0",x"70",x"05",x"38",x"20",x"c0",x"38",x"40",x"f8",x"70",x"98",x"98",x"98",x"18",x"0c",x"30",x"89",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"72",x"40",x"20",x"40",x"0c",x"40",x"0c",x"0c",x"20",x"40",x"60",x"c0",x"38",x"38",x"40",x"c7",x"38",x"40",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"40",x"38",x"40",x"40",x"40",x"40",x"89",x"90",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"72",x"40",x"20",x"40",x"0c",x"40",x"0c",x"20",x"5f",x"40",x"40",x"5f",x"90",x"90",x"0c",x"8a",x"86",x"82",x"8a",x"86",x"82",x"ca",x"38",x"20",x"40",x"40",x"8a",x"06",x"20",x"30",x"5f",x"90",x"0c",x"60",x"45",x"70",x"60",x"90",x"70",x"89",x"05",x"40",x"fc",x"00",x"c1",x"38",x"82",x"c2",x"38",x"38",x"60",x"45",x"80",x"c1",x"38",x"c9",x"38",x"98",x"18",x"50",x"38",x"89",x"ff",x"04",x"fc",x"00",x"c2",x"38",x"c2",x"38",x"40",x"40",x"40",x"80",x"70",x"20",x"89",x"0c",x"38",x"5f",x"70",x"10",x"40",x"c8",x"38",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"89",x"86",x"73",x"20",x"c3",x"38",x"60",x"0c",x"88",x"00",x"60",x"98",x"18",x"50",x"38",x"72",x"60",x"42",x"80",x"89",x"70",x"38",x"c1",x"38",x"89",x"82",x"88",x"89",x"05",x"05",x"30",x"5f",x"90",x"90",x"0c",x"ce",x"38",x"20",x"40",x"20",x"40",x"50",x"38",x"5c",x"90",x"90",x"90",x"0c",x"20",x"70",x"0c",x"89",x"90",x"ff",x"04",x"40",x"40",x"8f",x"7f",x"20",x"90",x"90",x"90",x"80",x"ef",x"c1",x"38",x"40",x"ef",x"c0",x"38",x"40",x"ff",x"7f",x"70",x"84",x"c0",x"38",x"70",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c1",x"38",x"60",x"85",x"c9",x"38",x"20",x"70",x"c0",x"38",x"70",x"60",x"c0",x"38",x"c0",x"38",x"04",x"c1",x"38",x"60",x"0c",x"c5",x"38",x"90",x"88",x"70",x"0c",x"40",x"0c",x"40",x"90",x"90",x"89",x"70",x"40",x"40",x"20",x"40",x"60",x"85",x"70",x"90",x"cc",x"38",x"40",x"70",x"70",x"40",x"20",x"40",x"8e",x"70",x"01",x"40",x"98",x"c9",x"38",x"40",x"70",x"98",x"01",x"90",x"70",x"40",x"40",x"98",x"98",x"70",x"01",x"98",x"01",x"8e",x"f0",x"81",x"90",x"70",x"20",x"40",x"04",x"40",x"40",x"98",x"00",x"40",x"42",x"50",x"38",x"60",x"86",x"05",x"c6",x"38",x"40",x"20",x"c6",x"38",x"38",x"20",x"40",x"20",x"0e",x"98",x"0c",x"40",x"45",x"44",x"60",x"43",x"45",x"90",x"8f",x"7f",x"40",x"05",x"40",x"98",x"06",x"60",x"41",x"85",x"60",x"42",x"f0",x"70",x"05",x"40",x"f8",x"70",x"ca",x"38",x"90",x"90",x"82",x"70",x"90",x"cb",x"38",x"c8",x"38",x"40",x"20",x"c0",x"38",x"40",x"85",x"60",x"41",x"c6",x"38",x"8f",x"6f",x"47",x"60",x"42",x"89",x"90",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"89",x"c6",x"38",x"0c",x"0c",x"40",x"74",x"40",x"90",x"82",x"0c",x"40",x"40",x"05",x"c0",x"38",x"90",x"98",x"98",x"98",x"0c",x"cd",x"38",x"40",x"05",x"40",x"40",x"40",x"05",x"90",x"0c",x"40",x"98",x"0c",x"70",x"80",x"60",x"47",x"70",x"40",x"c0",x"38",x"c0",x"38",x"98",x"05",x"05",x"20",x"20",x"70",x"06",x"60",x"41",x"70",x"04",x"01",x"38",x"40",x"70",x"98",x"98",x"98",x"18",x"53",x"38",x"40",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"89",x"85",x"80",x"0c",x"cb",x"38",x"40",x"70",x"82",x"8f",x"6f",x"4a",x"47",x"98",x"60",x"42",x"89",x"90",x"05",x"40",x"89",x"05",x"40",x"89",x"05",x"06",x"60",x"89",x"04",x"20",x"60",x"84",x"89",x"04",x"89",x"00",x"60",x"04",x"60",x"8b",x"89",x"47",x"90",x"90",x"c8",x"38",x"40",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"7f",x"d5",x"75",x"40",x"82",x"b3",x"73",x"20",x"40",x"00",x"40",x"8f",x"70",x"81",x"70",x"20",x"89",x"85",x"80",x"0c",x"c9",x"38",x"40",x"40",x"82",x"90",x"cf",x"38",x"5f",x"40",x"40",x"20",x"8b",x"00",x"60",x"84",x"84",x"18",x"20",x"20",x"40",x"8b",x"8b",x"84",x"80",x"04",x"88",x"00",x"89",x"89",x"00",x"00",x"30",x"5f",x"70",x"10",x"40",x"ce",x"38",x"40",x"50",x"38",x"70",x"c2",x"38",x"c1",x"38",x"40",x"89",x"05",x"40",x"89",x"05",x"40",x"20",x"40",x"89",x"05",x"40",x"7f",x"20",x"60",x"89",x"04",x"20",x"40",x"89",x"05",x"60",x"06",x"20",x"40",x"89",x"04",x"82",x"89",x"00",x"20",x"40",x"00",x"40",x"8f",x"70",x"04",x"60",x"8b",x"8b",x"89",x"89",x"82",x"61",x"47",x"c0",x"38",x"38",x"70",x"20",x"60",x"20",x"42",x"89",x"70",x"40",x"89",x"88",x"88",x"5f",x"05",x"82",x"8a",x"84",x"84",x"82",x"cd",x"38",x"40",x"20",x"30",x"5f",x"90",x"90",x"0c",x"cb",x"38",x"20",x"40",x"20",x"40",x"50",x"38",x"d4",x"6a",x"e3",x"11",x"1f",x"5e",x"e5",x"8d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"53",x"69",x"65",x"53",x"6b",x"20",x"66",x"61",x"20",x"20",x"61",x"65",x"66",x"63",x"6d",x"2e",x"6b",x"6c",x"74",x"20",x"20",x"61",x"65",x"66",x"63",x"6d",x"2e",x"72",x"6c",x"65",x"61",x"6e",x"6e",x"72",x"74",x"20",x"20",x"65",x"6b",x"32",x"65",x"72",x"63",x"75",x"61",x"65",x"73",x"72",x"72",x"72",x"00",x"76",x"64",x"6f",x"75",x"61",x"65",x"73",x"72",x"72",x"72",x"00",x"5d",x"4f",x"6c",x"20",x"20",x"30",x"2d",x"6f",x"20",x"30",x"34",x"5b",x"45",x"52",x"61",x"78",x"63",x"25",x"20",x"68",x"64",x"20",x"30",x"00",x"5d",x"4f",x"73",x"65",x"63",x"25",x"20",x"68",x"64",x"20",x"30",x"00",x"65",x"6b",x"7a",x"20",x"25",x"00",x"61",x"69",x"20",x"20",x"25",x"00",x"61",x"69",x"28",x"73",x"25",x"49",x"61",x"6e",x"65",x"20",x"66",x"52",x"21",x"73",x"78",x"74",x"6f",x"74",x"61",x"31",x"65",x"66",x"61",x"6c",x"72",x"6c",x"00",x"72",x"6f",x"20",x"20",x"25",x"00",x"70",x"72",x"72",x"6e",x"25",x"47",x"2e",x"20",x"70",x"62",x"43",x"67",x"33",x"61",x"52",x"41",x"33",x"69",x"29",x"6d",x"65",x"6c",x"20",x"20",x"00",x"6f",x"6c",x"74",x"20",x"25",x"53",x"4b",x"65",x"63",x"20",x"20",x"20",x"30",x"00",x"5d",x"6c",x"20",x"20",x"20",x"30",x"00",x"5d",x"6d",x"69",x"20",x"20",x"30",x"00",x"5d",x"73",x"65",x"20",x"20",x"30",x"00",x"5d",x"66",x"6c",x"20",x"20",x"30",x"00",x"72",x"20",x"72",x"6f",x"61",x"61",x"2e",x"65",x"61",x"2e",x"20",x"20",x"20",x"20",x"6f",x"6e",x"75",x"2e",x"6f",x"61",x"31",x"3a",x"20",x"73",x"00",x"25",x"72",x"73",x"74",x"65",x"43",x"6f",x"61",x"61",x"6f",x"61",x"6e",x"72",x"65",x"73",x"20",x"75",x"20",x"61",x"63",x"61",x"77",x"20",x"75",x"20",x"61",x"6f",x"70",x"66",x"2e",x"30",x"2d",x"2d",x"2b",x"00",x"2e",x"7a",x"2e",x"54",x"2e",x"65",x"2d",x"33",x"00",x"65",x"32",x"2e",x"31",x"35",x"34",x"2e",x"34",x"00",x"30",x"30",x"2e",x"30",x"30",x"31",x"00",x"34",x"32",x"4e",x"3e",x"32",x"36",x"61",x"65",x"69",x"6d",x"71",x"75",x"79",x"31",x"35",x"39",x"44",x"48",x"4c",x"50",x"54",x"58",x"00",x"00",x"00",x"00",x"90",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
signal rwea: std_logic_vector(3 downto 0);
signal rweb: std_logic_vector(3 downto 0);
signal memaread0: std_logic_vector(7 downto 0);
signal membread0: std_logic_vector(7 downto 0);
signal memaread1: std_logic_vector(7 downto 0);
signal membread1: std_logic_vector(7 downto 0);
signal memaread2: std_logic_vector(7 downto 0);
signal membread2: std_logic_vector(7 downto 0);
signal memaread3: std_logic_vector(7 downto 0);
signal membread3: std_logic_vector(7 downto 0);

begin
  rwea(0) <= WEA and MASKA(0);
  rweb(0) <= WEB and MASKB(0);
  rwea(1) <= WEA and MASKA(1);
  rweb(1) <= WEB and MASKB(1);
  rwea(2) <= WEA and MASKA(2);
  rweb(2) <= WEB and MASKB(2);
  rwea(3) <= WEA and MASKA(3);
  rweb(3) <= WEB and MASKB(3);
DOA(7 downto 0) <= memaread0;
DOB(7 downto 0) <= membread0;
DOA(15 downto 8) <= memaread1;
DOB(15 downto 8) <= membread1;
DOA(23 downto 16) <= memaread2;
DOB(23 downto 16) <= membread2;
DOA(31 downto 24) <= memaread3;
DOB(31 downto 24) <= membread3;

  process (clka)
  begin
    if rising_edge(clka) then
    if ENA='1' then
    if rwea(0)='1' then
      RAM0( conv_integer(ADDRA) ) := DIA(7 downto 0);
      end if;
    memaread0 <= RAM0(conv_integer(ADDRA)) ;
    end if;
    end if;
  end process;  

  process (clkb)
  begin
    if rising_edge(clkb) then
    if ENB='1' then
      if rweb(0)='1' then
         RAM0( conv_integer(ADDRB) ) := DIB(7 downto 0);
      end if;
      membread0 <= RAM0(conv_integer(ADDRB)) ;
    end if;
    end if;
  end process;  

  process (clka)
  begin
    if rising_edge(clka) then
    if ENA='1' then
    if rwea(1)='1' then
      RAM1( conv_integer(ADDRA) ) := DIA(15 downto 8);
      end if;
    memaread1 <= RAM1(conv_integer(ADDRA)) ;
    end if;
    end if;
  end process;  

  process (clkb)
  begin
    if rising_edge(clkb) then
    if ENB='1' then
      if rweb(1)='1' then
         RAM1( conv_integer(ADDRB) ) := DIB(15 downto 8);
      end if;
      membread1 <= RAM1(conv_integer(ADDRB)) ;
    end if;
    end if;
  end process;  

  process (clka)
  begin
    if rising_edge(clka) then
    if ENA='1' then
    if rwea(2)='1' then
      RAM2( conv_integer(ADDRA) ) := DIA(23 downto 16);
      end if;
    memaread2 <= RAM2(conv_integer(ADDRA)) ;
    end if;
    end if;
  end process;  

  process (clkb)
  begin
    if rising_edge(clkb) then
    if ENB='1' then
      if rweb(2)='1' then
         RAM2( conv_integer(ADDRB) ) := DIB(23 downto 16);
      end if;
      membread2 <= RAM2(conv_integer(ADDRB)) ;
    end if;
    end if;
  end process;  

  process (clka)
  begin
    if rising_edge(clka) then
    if ENA='1' then
    if rwea(3)='1' then
      RAM3( conv_integer(ADDRA) ) := DIA(31 downto 24);
      end if;
    memaread3 <= RAM3(conv_integer(ADDRA)) ;
    end if;
    end if;
  end process;  

  process (clkb)
  begin
    if rising_edge(clkb) then
    if ENB='1' then
      if rweb(3)='1' then
         RAM3( conv_integer(ADDRB) ) := DIB(31 downto 24);
      end if;
      membread3 <= RAM3(conv_integer(ADDRB)) ;
    end if;
    end if;
  end process;  
end behave;
